<!DOCTYPE html>
<!--[if IE]><![endif]-->
<html>
  
  <head>
    <meta charset="utf-8">
    <meta http-equiv="X-UA-Compatible" content="IE=edge,chrome=1">
    <title>Class MemberSuggestionsChangePolicyDetails
   </title>
    <meta name="viewport" content="width=device-width">
    <meta name="title" content="Class MemberSuggestionsChangePolicyDetails
   ">
    <meta name="generator" content="docfx 2.58.4.0">
    
    <link rel="shortcut icon" href="../../../favicon.ico">
    <link rel="stylesheet" href="../../../styles/docfx.vendor.css">
    <link rel="stylesheet" href="../../../styles/docfx.css">
    <link rel="stylesheet" href="../../../styles/main.css">
    <meta property="docfx:navrel" content="../../../toc.html">
    <meta property="docfx:tocrel" content="toc.html">
    
    
    
  </head>
  <body data-spy="scroll" data-target="#affix" data-offset="120">
    <div id="wrapper">
      <header>
        
        <nav id="autocollapse" class="navbar navbar-inverse ng-scope" role="navigation">
          <div class="container">
            <div class="navbar-header">
              <button type="button" class="navbar-toggle" data-toggle="collapse" data-target="#navbar">
                <span class="sr-only">Toggle navigation</span>
                <span class="icon-bar"></span>
                <span class="icon-bar"></span>
                <span class="icon-bar"></span>
              </button>
              
              <a class="navbar-brand" href="../../../index.html">
                <img id="logo" class="svg" src="../../../logo.svg" alt="">
              </a>
            </div>
            <div class="collapse navbar-collapse" id="navbar">
              <form class="navbar-form navbar-right" role="search" id="search">
                <div class="form-group">
                  <input type="text" class="form-control" id="search-query" placeholder="Search" autocomplete="off">
                </div>
              </form>
            </div>
          </div>
        </nav>
        
        <div class="subnav navbar navbar-default">
          <div class="container hide-when-search" id="breadcrumb">
            <ul class="breadcrumb">
              <li></li>
            </ul>
          </div>
        </div>
      </header>
      <div role="main" class="container body-content hide-when-search">
        
        <div class="sidenav hide-when-search">
          <a class="btn toc-toggle collapse" data-toggle="collapse" href="#sidetoggle" aria-expanded="false" aria-controls="sidetoggle">Show / Hide Table of Contents</a>
          <div class="sidetoggle collapse" id="sidetoggle">
            <div id="sidetoc"></div>
          </div>
        </div>
        <div class="article row grid-right">
          <div class="col-md-10">
            <article class="content wrap" id="_content" data-uid="Dropbox.Api.TeamLog.MemberSuggestionsChangePolicyDetails">
  
  
  <h1 id="Dropbox_Api_TeamLog_MemberSuggestionsChangePolicyDetails" data-uid="Dropbox.Api.TeamLog.MemberSuggestionsChangePolicyDetails" class="text-break">Class MemberSuggestionsChangePolicyDetails
  </h1>
  <div class="markdown level0 summary"><p>Enabled/disabled option for team members to suggest people to add to team.</p>
</div>
  <div class="markdown level0 conceptual"></div>
  <div class="inheritance">
    <h5>Inheritance</h5>
    <div class="level0"><span class="xref">System.Object</span></div>
    <div class="level1"><span class="xref">MemberSuggestionsChangePolicyDetails</span></div>
  </div>
  <div class="inheritedMembers">
    <h5>Inherited Members</h5>
    <div>
      <span class="xref">System.Object.Equals(System.Object)</span>
    </div>
    <div>
      <span class="xref">System.Object.Equals(System.Object, System.Object)</span>
    </div>
    <div>
      <span class="xref">System.Object.GetHashCode()</span>
    </div>
    <div>
      <span class="xref">System.Object.GetType()</span>
    </div>
    <div>
      <span class="xref">System.Object.MemberwiseClone()</span>
    </div>
    <div>
      <span class="xref">System.Object.ReferenceEquals(System.Object, System.Object)</span>
    </div>
    <div>
      <span class="xref">System.Object.ToString()</span>
    </div>
  </div>
  <h6><strong>Namespace</strong>: <a class="xref" href="Dropbox.Api.TeamLog.html">Dropbox.Api.TeamLog</a></h6>
  <h6><strong>Assembly</strong>: Dropbox.Api.dll</h6>
  <h5 id="Dropbox_Api_TeamLog_MemberSuggestionsChangePolicyDetails_syntax">Syntax</h5>
  <div class="codewrapper">
    <pre><code class="lang-csharp hljs">public class MemberSuggestionsChangePolicyDetails</code></pre>
  </div>
  <h3 id="constructors">Constructors
  </h3>
  <span class="small pull-right mobile-hide">
    <span class="divider">|</span>
    <a href="https://github.com/dropbox/dropbox-sdk-dotnet/new/doc_fx_integration/apiSpec/new?filename=Dropbox_Api_TeamLog_MemberSuggestionsChangePolicyDetails__ctor_Dropbox_Api_TeamLog_MemberSuggestionsPolicy_Dropbox_Api_TeamLog_MemberSuggestionsPolicy_.md&amp;value=---%0Auid%3A%20Dropbox.Api.TeamLog.MemberSuggestionsChangePolicyDetails.%23ctor(Dropbox.Api.TeamLog.MemberSuggestionsPolicy%2CDropbox.Api.TeamLog.MemberSuggestionsPolicy)%0Asummary%3A%20'*You%20can%20override%20summary%20for%20the%20API%20here%20using%20*MARKDOWN*%20syntax'%0A---%0A%0A*Please%20type%20below%20more%20information%20about%20this%20API%3A*%0A%0A">Improve this Doc</a>
  </span>
  <span class="small pull-right mobile-hide">
    <a href="https://github.com/dropbox/dropbox-sdk-dotnet/blob/doc_fx_integration/dropbox-sdk-dotnet/Dropbox.Api/Generated/TeamLog/MemberSuggestionsChangePolicyDetails.cs/#L37">View Source</a>
  </span>
  <a id="Dropbox_Api_TeamLog_MemberSuggestionsChangePolicyDetails__ctor_" data-uid="Dropbox.Api.TeamLog.MemberSuggestionsChangePolicyDetails.#ctor*"></a>
  <h4 id="Dropbox_Api_TeamLog_MemberSuggestionsChangePolicyDetails__ctor_Dropbox_Api_TeamLog_MemberSuggestionsPolicy_Dropbox_Api_TeamLog_MemberSuggestionsPolicy_" data-uid="Dropbox.Api.TeamLog.MemberSuggestionsChangePolicyDetails.#ctor(Dropbox.Api.TeamLog.MemberSuggestionsPolicy,Dropbox.Api.TeamLog.MemberSuggestionsPolicy)">MemberSuggestionsChangePolicyDetails(MemberSuggestionsPolicy, MemberSuggestionsPolicy)</h4>
  <div class="markdown level1 summary"><p>Initializes a new instance of the <a class="xref" href="Dropbox.Api.TeamLog.MemberSuggestionsChangePolicyDetails.html">MemberSuggestionsChangePolicyDetails</a> class.</p>
</div>
  <div class="markdown level1 conceptual"></div>
  <h5 class="decalaration">Declaration</h5>
  <div class="codewrapper">
    <pre><code class="lang-csharp hljs">public MemberSuggestionsChangePolicyDetails(MemberSuggestionsPolicy newValue, MemberSuggestionsPolicy previousValue = null)</code></pre>
  </div>
  <h5 class="parameters">Parameters</h5>
  <table class="table table-bordered table-striped table-condensed">
    <thead>
      <tr>
        <th>Type</th>
        <th>Name</th>
        <th>Description</th>
      </tr>
    </thead>
    <tbody>
      <tr>
        <td><a class="xref" href="Dropbox.Api.TeamLog.MemberSuggestionsPolicy.html">MemberSuggestionsPolicy</a></td>
        <td><span class="parametername">newValue</span></td>
        <td><p sourcefile="gh-pages/obj/api/Dropbox.Api.TeamLog.MemberSuggestionsChangePolicyDetails.yml" sourcestartlinenumber="1" sourceendlinenumber="1">New team member suggestions policy.</p>
</td>
      </tr>
      <tr>
        <td><a class="xref" href="Dropbox.Api.TeamLog.MemberSuggestionsPolicy.html">MemberSuggestionsPolicy</a></td>
        <td><span class="parametername">previousValue</span></td>
        <td><p sourcefile="gh-pages/obj/api/Dropbox.Api.TeamLog.MemberSuggestionsChangePolicyDetails.yml" sourcestartlinenumber="1" sourceendlinenumber="2">Previous team member suggestions policy. Might be
missing due to historical data gap.</p>
</td>
      </tr>
    </tbody>
  </table>
  <h3 id="properties">Properties
  </h3>
  <span class="small pull-right mobile-hide">
    <span class="divider">|</span>
    <a href="https://github.com/dropbox/dropbox-sdk-dotnet/new/doc_fx_integration/apiSpec/new?filename=Dropbox_Api_TeamLog_MemberSuggestionsChangePolicyDetails_NewValue.md&amp;value=---%0Auid%3A%20Dropbox.Api.TeamLog.MemberSuggestionsChangePolicyDetails.NewValue%0Asummary%3A%20'*You%20can%20override%20summary%20for%20the%20API%20here%20using%20*MARKDOWN*%20syntax'%0A---%0A%0A*Please%20type%20below%20more%20information%20about%20this%20API%3A*%0A%0A">Improve this Doc</a>
  </span>
  <span class="small pull-right mobile-hide">
    <a href="https://github.com/dropbox/dropbox-sdk-dotnet/blob/doc_fx_integration/dropbox-sdk-dotnet/Dropbox.Api/Generated/TeamLog/MemberSuggestionsChangePolicyDetails.cs/#L63">View Source</a>
  </span>
  <a id="Dropbox_Api_TeamLog_MemberSuggestionsChangePolicyDetails_NewValue_" data-uid="Dropbox.Api.TeamLog.MemberSuggestionsChangePolicyDetails.NewValue*"></a>
  <h4 id="Dropbox_Api_TeamLog_MemberSuggestionsChangePolicyDetails_NewValue" data-uid="Dropbox.Api.TeamLog.MemberSuggestionsChangePolicyDetails.NewValue">NewValue</h4>
  <div class="markdown level1 summary"><p>New team member suggestions policy.</p>
</div>
  <div class="markdown level1 conceptual"></div>
  <h5 class="decalaration">Declaration</h5>
  <div class="codewrapper">
    <pre><code class="lang-csharp hljs">public MemberSuggestionsPolicy NewValue { get; protected set; }</code></pre>
  </div>
  <h5 class="propertyValue">Property Value</h5>
  <table class="table table-bordered table-striped table-condensed">
    <thead>
      <tr>
        <th>Type</th>
        <th>Description</th>
      </tr>
    </thead>
    <tbody>
      <tr>
        <td><a class="xref" href="Dropbox.Api.TeamLog.MemberSuggestionsPolicy.html">MemberSuggestionsPolicy</a></td>
        <td></td>
      </tr>
    </tbody>
  </table>
  <span class="small pull-right mobile-hide">
    <span class="divider">|</span>
    <a href="https://github.com/dropbox/dropbox-sdk-dotnet/new/doc_fx_integration/apiSpec/new?filename=Dropbox_Api_TeamLog_MemberSuggestionsChangePolicyDetails_PreviousValue.md&amp;value=---%0Auid%3A%20Dropbox.Api.TeamLog.MemberSuggestionsChangePolicyDetails.PreviousValue%0Asummary%3A%20'*You%20can%20override%20summary%20for%20the%20API%20here%20using%20*MARKDOWN*%20syntax'%0A---%0A%0A*Please%20type%20below%20more%20information%20about%20this%20API%3A*%0A%0A">Improve this Doc</a>
  </span>
  <span class="small pull-right mobile-hide">
    <a href="https://github.com/dropbox/dropbox-sdk-dotnet/blob/doc_fx_integration/dropbox-sdk-dotnet/Dropbox.Api/Generated/TeamLog/MemberSuggestionsChangePolicyDetails.cs/#L69">View Source</a>
  </span>
  <a id="Dropbox_Api_TeamLog_MemberSuggestionsChangePolicyDetails_PreviousValue_" data-uid="Dropbox.Api.TeamLog.MemberSuggestionsChangePolicyDetails.PreviousValue*"></a>
  <h4 id="Dropbox_Api_TeamLog_MemberSuggestionsChangePolicyDetails_PreviousValue" data-uid="Dropbox.Api.TeamLog.MemberSuggestionsChangePolicyDetails.PreviousValue">PreviousValue</h4>
  <div class="markdown level1 summary"><p>Previous team member suggestions policy. Might be missing due to historical
data gap.</p>
</div>
  <div class="markdown level1 conceptual"></div>
  <h5 class="decalaration">Declaration</h5>
  <div class="codewrapper">
    <pre><code class="lang-csharp hljs">public MemberSuggestionsPolicy PreviousValue { get; protected set; }</code></pre>
  </div>
  <h5 class="propertyValue">Property Value</h5>
  <table class="table table-bordered table-striped table-condensed">
    <thead>
      <tr>
        <th>Type</th>
        <th>Description</th>
      </tr>
    </thead>
    <tbody>
      <tr>
        <td><a class="xref" href="Dropbox.Api.TeamLog.MemberSuggestionsPolicy.html">MemberSuggestionsPolicy</a></td>
        <td></td>
      </tr>
    </tbody>
  </table>
</article>
          </div>
          
          <div class="hidden-sm col-md-2" role="complementary">
            <div class="sideaffix">
              <div class="contribution">
                <ul class="nav">
                  <li>
                    <a href="https://github.com/dropbox/dropbox-sdk-dotnet/new/doc_fx_integration/apiSpec/new?filename=Dropbox_Api_TeamLog_MemberSuggestionsChangePolicyDetails.md&amp;value=---%0Auid%3A%20Dropbox.Api.TeamLog.MemberSuggestionsChangePolicyDetails%0Asummary%3A%20'*You%20can%20override%20summary%20for%20the%20API%20here%20using%20*MARKDOWN*%20syntax'%0A---%0A%0A*Please%20type%20below%20more%20information%20about%20this%20API%3A*%0A%0A" class="contribution-link">Improve this Doc</a>
                  </li>
                  <li>
                    <a href="https://github.com/dropbox/dropbox-sdk-dotnet/blob/doc_fx_integration/dropbox-sdk-dotnet/Dropbox.Api/Generated/TeamLog/MemberSuggestionsChangePolicyDetails.cs/#L16" class="contribution-link">View Source</a>
                  </li>
                </ul>
              </div>
              <nav class="bs-docs-sidebar hidden-print hidden-xs hidden-sm affix" id="affix">
                <h5>In This Article</h5>
                <div></div>
              </nav>
            </div>
          </div>
        </div>
      </div>
      
      <footer>
        <div class="grad-bottom"></div>
        <div class="footer">
          <div class="container">
            <span class="pull-right">
              <a href="#top">Back to top</a>
            </span>
            
            <span>Generated by <strong>DocFX</strong></span>
          </div>
        </div>
      </footer>
    </div>
    
    <script type="text/javascript" src="../../../styles/docfx.vendor.js"></script>
    <script type="text/javascript" src="../../../styles/docfx.js"></script>
    <script type="text/javascript" src="../../../styles/main.js"></script>
  </body>
</html>
