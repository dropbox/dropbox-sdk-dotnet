﻿<!DOCTYPE html>
<!--[if IE]><![endif]-->
<html>
  
  <head>
    <meta charset="utf-8">
    <meta http-equiv="X-UA-Compatible" content="IE=edge,chrome=1">
    <title>Class EventTypeArg.SharedLinkRemoveExpiry
   </title>
    <meta name="viewport" content="width=device-width">
    <meta name="title" content="Class EventTypeArg.SharedLinkRemoveExpiry
   ">
    <meta name="generator" content="docfx 2.58.4.0">
    
    <link rel="shortcut icon" href="../../../favicon.ico">
    <link rel="stylesheet" href="../../../styles/docfx.vendor.css">
    <link rel="stylesheet" href="../../../styles/docfx.css">
    <link rel="stylesheet" href="../../../styles/main.css">
    <meta property="docfx:navrel" content="../../../toc.html">
    <meta property="docfx:tocrel" content="toc.html">
    
    
    
  </head>
  <body data-spy="scroll" data-target="#affix" data-offset="120">
    <div id="wrapper">
      <header>
        
        <nav id="autocollapse" class="navbar navbar-inverse ng-scope" role="navigation">
          <div class="container">
            <div class="navbar-header">
              <button type="button" class="navbar-toggle" data-toggle="collapse" data-target="#navbar">
                <span class="sr-only">Toggle navigation</span>
                <span class="icon-bar"></span>
                <span class="icon-bar"></span>
                <span class="icon-bar"></span>
              </button>
              
              <a class="navbar-brand" href="../../../index.html">
                <img id="logo" class="svg" src="../../../logo.svg" alt="">
              </a>
            </div>
            <div class="collapse navbar-collapse" id="navbar">
              <form class="navbar-form navbar-right" role="search" id="search">
                <div class="form-group">
                  <input type="text" class="form-control" id="search-query" placeholder="Search" autocomplete="off">
                </div>
              </form>
            </div>
          </div>
        </nav>
        
        <div class="subnav navbar navbar-default">
          <div class="container hide-when-search" id="breadcrumb">
            <ul class="breadcrumb">
              <li></li>
            </ul>
          </div>
        </div>
      </header>
      <div role="main" class="container body-content hide-when-search">
        
        <div class="sidenav hide-when-search">
          <a class="btn toc-toggle collapse" data-toggle="collapse" href="#sidetoggle" aria-expanded="false" aria-controls="sidetoggle">Show / Hide Table of Contents</a>
          <div class="sidetoggle collapse" id="sidetoggle">
            <div id="sidetoc"></div>
          </div>
        </div>
        <div class="article row grid-right">
          <div class="col-md-10">
            <article class="content wrap" id="_content" data-uid="Dropbox.Api.TeamLog.EventTypeArg.SharedLinkRemoveExpiry">
  
  
  <h1 id="Dropbox_Api_TeamLog_EventTypeArg_SharedLinkRemoveExpiry" data-uid="Dropbox.Api.TeamLog.EventTypeArg.SharedLinkRemoveExpiry" class="text-break">Class EventTypeArg.SharedLinkRemoveExpiry
  </h1>
  <div class="markdown level0 summary"><p>(sharing) Removed shared link expiration date</p>
</div>
  <div class="markdown level0 conceptual"></div>
  <div class="inheritance">
    <h5>Inheritance</h5>
    <div class="level0"><span class="xref">System.Object</span></div>
    <div class="level1"><a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html">EventTypeArg</a></div>
    <div class="level2"><span class="xref">EventTypeArg.SharedLinkRemoveExpiry</span></div>
  </div>
  <div class="inheritedMembers">
    <h5>Inherited Members</h5>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsAdminAlertingAlertStateChanged">EventTypeArg.IsAdminAlertingAlertStateChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsAdminAlertingAlertStateChanged">EventTypeArg.AsAdminAlertingAlertStateChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsAdminAlertingChangedAlertConfig">EventTypeArg.IsAdminAlertingChangedAlertConfig</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsAdminAlertingChangedAlertConfig">EventTypeArg.AsAdminAlertingChangedAlertConfig</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsAdminAlertingTriggeredAlert">EventTypeArg.IsAdminAlertingTriggeredAlert</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsAdminAlertingTriggeredAlert">EventTypeArg.AsAdminAlertingTriggeredAlert</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsAppBlockedByPermissions">EventTypeArg.IsAppBlockedByPermissions</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsAppBlockedByPermissions">EventTypeArg.AsAppBlockedByPermissions</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsAppLinkTeam">EventTypeArg.IsAppLinkTeam</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsAppLinkTeam">EventTypeArg.AsAppLinkTeam</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsAppLinkUser">EventTypeArg.IsAppLinkUser</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsAppLinkUser">EventTypeArg.AsAppLinkUser</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsAppUnlinkTeam">EventTypeArg.IsAppUnlinkTeam</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsAppUnlinkTeam">EventTypeArg.AsAppUnlinkTeam</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsAppUnlinkUser">EventTypeArg.IsAppUnlinkUser</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsAppUnlinkUser">EventTypeArg.AsAppUnlinkUser</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsIntegrationConnected">EventTypeArg.IsIntegrationConnected</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsIntegrationConnected">EventTypeArg.AsIntegrationConnected</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsIntegrationDisconnected">EventTypeArg.IsIntegrationDisconnected</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsIntegrationDisconnected">EventTypeArg.AsIntegrationDisconnected</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileAddComment">EventTypeArg.IsFileAddComment</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileAddComment">EventTypeArg.AsFileAddComment</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileChangeCommentSubscription">EventTypeArg.IsFileChangeCommentSubscription</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileChangeCommentSubscription">EventTypeArg.AsFileChangeCommentSubscription</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileDeleteComment">EventTypeArg.IsFileDeleteComment</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileDeleteComment">EventTypeArg.AsFileDeleteComment</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileEditComment">EventTypeArg.IsFileEditComment</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileEditComment">EventTypeArg.AsFileEditComment</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileLikeComment">EventTypeArg.IsFileLikeComment</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileLikeComment">EventTypeArg.AsFileLikeComment</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileResolveComment">EventTypeArg.IsFileResolveComment</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileResolveComment">EventTypeArg.AsFileResolveComment</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileUnlikeComment">EventTypeArg.IsFileUnlikeComment</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileUnlikeComment">EventTypeArg.AsFileUnlikeComment</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileUnresolveComment">EventTypeArg.IsFileUnresolveComment</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileUnresolveComment">EventTypeArg.AsFileUnresolveComment</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsGovernancePolicyAddFolders">EventTypeArg.IsGovernancePolicyAddFolders</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsGovernancePolicyAddFolders">EventTypeArg.AsGovernancePolicyAddFolders</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsGovernancePolicyAddFolderFailed">EventTypeArg.IsGovernancePolicyAddFolderFailed</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsGovernancePolicyAddFolderFailed">EventTypeArg.AsGovernancePolicyAddFolderFailed</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsGovernancePolicyContentDisposed">EventTypeArg.IsGovernancePolicyContentDisposed</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsGovernancePolicyContentDisposed">EventTypeArg.AsGovernancePolicyContentDisposed</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsGovernancePolicyCreate">EventTypeArg.IsGovernancePolicyCreate</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsGovernancePolicyCreate">EventTypeArg.AsGovernancePolicyCreate</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsGovernancePolicyDelete">EventTypeArg.IsGovernancePolicyDelete</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsGovernancePolicyDelete">EventTypeArg.AsGovernancePolicyDelete</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsGovernancePolicyEditDetails">EventTypeArg.IsGovernancePolicyEditDetails</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsGovernancePolicyEditDetails">EventTypeArg.AsGovernancePolicyEditDetails</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsGovernancePolicyEditDuration">EventTypeArg.IsGovernancePolicyEditDuration</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsGovernancePolicyEditDuration">EventTypeArg.AsGovernancePolicyEditDuration</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsGovernancePolicyExportCreated">EventTypeArg.IsGovernancePolicyExportCreated</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsGovernancePolicyExportCreated">EventTypeArg.AsGovernancePolicyExportCreated</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsGovernancePolicyExportRemoved">EventTypeArg.IsGovernancePolicyExportRemoved</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsGovernancePolicyExportRemoved">EventTypeArg.AsGovernancePolicyExportRemoved</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsGovernancePolicyRemoveFolders">EventTypeArg.IsGovernancePolicyRemoveFolders</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsGovernancePolicyRemoveFolders">EventTypeArg.AsGovernancePolicyRemoveFolders</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsGovernancePolicyReportCreated">EventTypeArg.IsGovernancePolicyReportCreated</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsGovernancePolicyReportCreated">EventTypeArg.AsGovernancePolicyReportCreated</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsGovernancePolicyZipPartDownloaded">EventTypeArg.IsGovernancePolicyZipPartDownloaded</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsGovernancePolicyZipPartDownloaded">EventTypeArg.AsGovernancePolicyZipPartDownloaded</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsLegalHoldsActivateAHold">EventTypeArg.IsLegalHoldsActivateAHold</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsLegalHoldsActivateAHold">EventTypeArg.AsLegalHoldsActivateAHold</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsLegalHoldsAddMembers">EventTypeArg.IsLegalHoldsAddMembers</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsLegalHoldsAddMembers">EventTypeArg.AsLegalHoldsAddMembers</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsLegalHoldsChangeHoldDetails">EventTypeArg.IsLegalHoldsChangeHoldDetails</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsLegalHoldsChangeHoldDetails">EventTypeArg.AsLegalHoldsChangeHoldDetails</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsLegalHoldsChangeHoldName">EventTypeArg.IsLegalHoldsChangeHoldName</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsLegalHoldsChangeHoldName">EventTypeArg.AsLegalHoldsChangeHoldName</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsLegalHoldsExportAHold">EventTypeArg.IsLegalHoldsExportAHold</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsLegalHoldsExportAHold">EventTypeArg.AsLegalHoldsExportAHold</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsLegalHoldsExportCancelled">EventTypeArg.IsLegalHoldsExportCancelled</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsLegalHoldsExportCancelled">EventTypeArg.AsLegalHoldsExportCancelled</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsLegalHoldsExportDownloaded">EventTypeArg.IsLegalHoldsExportDownloaded</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsLegalHoldsExportDownloaded">EventTypeArg.AsLegalHoldsExportDownloaded</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsLegalHoldsExportRemoved">EventTypeArg.IsLegalHoldsExportRemoved</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsLegalHoldsExportRemoved">EventTypeArg.AsLegalHoldsExportRemoved</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsLegalHoldsReleaseAHold">EventTypeArg.IsLegalHoldsReleaseAHold</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsLegalHoldsReleaseAHold">EventTypeArg.AsLegalHoldsReleaseAHold</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsLegalHoldsRemoveMembers">EventTypeArg.IsLegalHoldsRemoveMembers</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsLegalHoldsRemoveMembers">EventTypeArg.AsLegalHoldsRemoveMembers</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsLegalHoldsReportAHold">EventTypeArg.IsLegalHoldsReportAHold</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsLegalHoldsReportAHold">EventTypeArg.AsLegalHoldsReportAHold</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDeviceChangeIpDesktop">EventTypeArg.IsDeviceChangeIpDesktop</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDeviceChangeIpDesktop">EventTypeArg.AsDeviceChangeIpDesktop</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDeviceChangeIpMobile">EventTypeArg.IsDeviceChangeIpMobile</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDeviceChangeIpMobile">EventTypeArg.AsDeviceChangeIpMobile</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDeviceChangeIpWeb">EventTypeArg.IsDeviceChangeIpWeb</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDeviceChangeIpWeb">EventTypeArg.AsDeviceChangeIpWeb</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDeviceDeleteOnUnlinkFail">EventTypeArg.IsDeviceDeleteOnUnlinkFail</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDeviceDeleteOnUnlinkFail">EventTypeArg.AsDeviceDeleteOnUnlinkFail</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDeviceDeleteOnUnlinkSuccess">EventTypeArg.IsDeviceDeleteOnUnlinkSuccess</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDeviceDeleteOnUnlinkSuccess">EventTypeArg.AsDeviceDeleteOnUnlinkSuccess</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDeviceLinkFail">EventTypeArg.IsDeviceLinkFail</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDeviceLinkFail">EventTypeArg.AsDeviceLinkFail</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDeviceLinkSuccess">EventTypeArg.IsDeviceLinkSuccess</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDeviceLinkSuccess">EventTypeArg.AsDeviceLinkSuccess</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDeviceManagementDisabled">EventTypeArg.IsDeviceManagementDisabled</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDeviceManagementDisabled">EventTypeArg.AsDeviceManagementDisabled</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDeviceManagementEnabled">EventTypeArg.IsDeviceManagementEnabled</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDeviceManagementEnabled">EventTypeArg.AsDeviceManagementEnabled</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDeviceSyncBackupStatusChanged">EventTypeArg.IsDeviceSyncBackupStatusChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDeviceSyncBackupStatusChanged">EventTypeArg.AsDeviceSyncBackupStatusChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDeviceUnlink">EventTypeArg.IsDeviceUnlink</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDeviceUnlink">EventTypeArg.AsDeviceUnlink</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDropboxPasswordsExported">EventTypeArg.IsDropboxPasswordsExported</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDropboxPasswordsExported">EventTypeArg.AsDropboxPasswordsExported</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDropboxPasswordsNewDeviceEnrolled">EventTypeArg.IsDropboxPasswordsNewDeviceEnrolled</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDropboxPasswordsNewDeviceEnrolled">EventTypeArg.AsDropboxPasswordsNewDeviceEnrolled</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsEmmRefreshAuthToken">EventTypeArg.IsEmmRefreshAuthToken</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsEmmRefreshAuthToken">EventTypeArg.AsEmmRefreshAuthToken</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsExternalDriveBackupEligibilityStatusChecked">EventTypeArg.IsExternalDriveBackupEligibilityStatusChecked</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsExternalDriveBackupEligibilityStatusChecked">EventTypeArg.AsExternalDriveBackupEligibilityStatusChecked</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsExternalDriveBackupStatusChanged">EventTypeArg.IsExternalDriveBackupStatusChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsExternalDriveBackupStatusChanged">EventTypeArg.AsExternalDriveBackupStatusChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsAccountCaptureChangeAvailability">EventTypeArg.IsAccountCaptureChangeAvailability</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsAccountCaptureChangeAvailability">EventTypeArg.AsAccountCaptureChangeAvailability</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsAccountCaptureMigrateAccount">EventTypeArg.IsAccountCaptureMigrateAccount</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsAccountCaptureMigrateAccount">EventTypeArg.AsAccountCaptureMigrateAccount</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsAccountCaptureNotificationEmailsSent">EventTypeArg.IsAccountCaptureNotificationEmailsSent</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsAccountCaptureNotificationEmailsSent">EventTypeArg.AsAccountCaptureNotificationEmailsSent</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsAccountCaptureRelinquishAccount">EventTypeArg.IsAccountCaptureRelinquishAccount</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsAccountCaptureRelinquishAccount">EventTypeArg.AsAccountCaptureRelinquishAccount</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDisabledDomainInvites">EventTypeArg.IsDisabledDomainInvites</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDisabledDomainInvites">EventTypeArg.AsDisabledDomainInvites</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDomainInvitesApproveRequestToJoinTeam">EventTypeArg.IsDomainInvitesApproveRequestToJoinTeam</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDomainInvitesApproveRequestToJoinTeam">EventTypeArg.AsDomainInvitesApproveRequestToJoinTeam</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDomainInvitesDeclineRequestToJoinTeam">EventTypeArg.IsDomainInvitesDeclineRequestToJoinTeam</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDomainInvitesDeclineRequestToJoinTeam">EventTypeArg.AsDomainInvitesDeclineRequestToJoinTeam</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDomainInvitesEmailExistingUsers">EventTypeArg.IsDomainInvitesEmailExistingUsers</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDomainInvitesEmailExistingUsers">EventTypeArg.AsDomainInvitesEmailExistingUsers</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDomainInvitesRequestToJoinTeam">EventTypeArg.IsDomainInvitesRequestToJoinTeam</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDomainInvitesRequestToJoinTeam">EventTypeArg.AsDomainInvitesRequestToJoinTeam</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDomainInvitesSetInviteNewUserPrefToNo">EventTypeArg.IsDomainInvitesSetInviteNewUserPrefToNo</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDomainInvitesSetInviteNewUserPrefToNo">EventTypeArg.AsDomainInvitesSetInviteNewUserPrefToNo</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDomainInvitesSetInviteNewUserPrefToYes">EventTypeArg.IsDomainInvitesSetInviteNewUserPrefToYes</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDomainInvitesSetInviteNewUserPrefToYes">EventTypeArg.AsDomainInvitesSetInviteNewUserPrefToYes</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDomainVerificationAddDomainFail">EventTypeArg.IsDomainVerificationAddDomainFail</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDomainVerificationAddDomainFail">EventTypeArg.AsDomainVerificationAddDomainFail</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDomainVerificationAddDomainSuccess">EventTypeArg.IsDomainVerificationAddDomainSuccess</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDomainVerificationAddDomainSuccess">EventTypeArg.AsDomainVerificationAddDomainSuccess</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDomainVerificationRemoveDomain">EventTypeArg.IsDomainVerificationRemoveDomain</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDomainVerificationRemoveDomain">EventTypeArg.AsDomainVerificationRemoveDomain</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsEnabledDomainInvites">EventTypeArg.IsEnabledDomainInvites</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsEnabledDomainInvites">EventTypeArg.AsEnabledDomainInvites</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsApplyNamingConvention">EventTypeArg.IsApplyNamingConvention</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsApplyNamingConvention">EventTypeArg.AsApplyNamingConvention</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsCreateFolder">EventTypeArg.IsCreateFolder</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsCreateFolder">EventTypeArg.AsCreateFolder</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileAdd">EventTypeArg.IsFileAdd</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileAdd">EventTypeArg.AsFileAdd</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileCopy">EventTypeArg.IsFileCopy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileCopy">EventTypeArg.AsFileCopy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileDelete">EventTypeArg.IsFileDelete</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileDelete">EventTypeArg.AsFileDelete</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileDownload">EventTypeArg.IsFileDownload</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileDownload">EventTypeArg.AsFileDownload</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileEdit">EventTypeArg.IsFileEdit</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileEdit">EventTypeArg.AsFileEdit</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileGetCopyReference">EventTypeArg.IsFileGetCopyReference</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileGetCopyReference">EventTypeArg.AsFileGetCopyReference</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileLockingLockStatusChanged">EventTypeArg.IsFileLockingLockStatusChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileLockingLockStatusChanged">EventTypeArg.AsFileLockingLockStatusChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileMove">EventTypeArg.IsFileMove</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileMove">EventTypeArg.AsFileMove</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFilePermanentlyDelete">EventTypeArg.IsFilePermanentlyDelete</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFilePermanentlyDelete">EventTypeArg.AsFilePermanentlyDelete</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFilePreview">EventTypeArg.IsFilePreview</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFilePreview">EventTypeArg.AsFilePreview</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileRename">EventTypeArg.IsFileRename</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileRename">EventTypeArg.AsFileRename</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileRestore">EventTypeArg.IsFileRestore</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileRestore">EventTypeArg.AsFileRestore</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileRevert">EventTypeArg.IsFileRevert</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileRevert">EventTypeArg.AsFileRevert</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileRollbackChanges">EventTypeArg.IsFileRollbackChanges</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileRollbackChanges">EventTypeArg.AsFileRollbackChanges</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileSaveCopyReference">EventTypeArg.IsFileSaveCopyReference</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileSaveCopyReference">EventTypeArg.AsFileSaveCopyReference</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFolderOverviewDescriptionChanged">EventTypeArg.IsFolderOverviewDescriptionChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFolderOverviewDescriptionChanged">EventTypeArg.AsFolderOverviewDescriptionChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFolderOverviewItemPinned">EventTypeArg.IsFolderOverviewItemPinned</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFolderOverviewItemPinned">EventTypeArg.AsFolderOverviewItemPinned</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFolderOverviewItemUnpinned">EventTypeArg.IsFolderOverviewItemUnpinned</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFolderOverviewItemUnpinned">EventTypeArg.AsFolderOverviewItemUnpinned</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsObjectLabelAdded">EventTypeArg.IsObjectLabelAdded</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsObjectLabelAdded">EventTypeArg.AsObjectLabelAdded</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsObjectLabelRemoved">EventTypeArg.IsObjectLabelRemoved</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsObjectLabelRemoved">EventTypeArg.AsObjectLabelRemoved</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsObjectLabelUpdatedValue">EventTypeArg.IsObjectLabelUpdatedValue</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsObjectLabelUpdatedValue">EventTypeArg.AsObjectLabelUpdatedValue</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsOrganizeFolderWithTidy">EventTypeArg.IsOrganizeFolderWithTidy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsOrganizeFolderWithTidy">EventTypeArg.AsOrganizeFolderWithTidy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsRewindFolder">EventTypeArg.IsRewindFolder</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsRewindFolder">EventTypeArg.AsRewindFolder</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsUndoNamingConvention">EventTypeArg.IsUndoNamingConvention</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsUndoNamingConvention">EventTypeArg.AsUndoNamingConvention</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsUndoOrganizeFolderWithTidy">EventTypeArg.IsUndoOrganizeFolderWithTidy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsUndoOrganizeFolderWithTidy">EventTypeArg.AsUndoOrganizeFolderWithTidy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsUserTagsAdded">EventTypeArg.IsUserTagsAdded</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsUserTagsAdded">EventTypeArg.AsUserTagsAdded</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsUserTagsRemoved">EventTypeArg.IsUserTagsRemoved</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsUserTagsRemoved">EventTypeArg.AsUserTagsRemoved</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsEmailIngestReceiveFile">EventTypeArg.IsEmailIngestReceiveFile</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsEmailIngestReceiveFile">EventTypeArg.AsEmailIngestReceiveFile</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileRequestChange">EventTypeArg.IsFileRequestChange</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileRequestChange">EventTypeArg.AsFileRequestChange</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileRequestClose">EventTypeArg.IsFileRequestClose</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileRequestClose">EventTypeArg.AsFileRequestClose</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileRequestCreate">EventTypeArg.IsFileRequestCreate</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileRequestCreate">EventTypeArg.AsFileRequestCreate</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileRequestDelete">EventTypeArg.IsFileRequestDelete</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileRequestDelete">EventTypeArg.AsFileRequestDelete</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileRequestReceiveFile">EventTypeArg.IsFileRequestReceiveFile</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileRequestReceiveFile">EventTypeArg.AsFileRequestReceiveFile</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsGroupAddExternalId">EventTypeArg.IsGroupAddExternalId</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsGroupAddExternalId">EventTypeArg.AsGroupAddExternalId</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsGroupAddMember">EventTypeArg.IsGroupAddMember</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsGroupAddMember">EventTypeArg.AsGroupAddMember</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsGroupChangeExternalId">EventTypeArg.IsGroupChangeExternalId</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsGroupChangeExternalId">EventTypeArg.AsGroupChangeExternalId</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsGroupChangeManagementType">EventTypeArg.IsGroupChangeManagementType</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsGroupChangeManagementType">EventTypeArg.AsGroupChangeManagementType</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsGroupChangeMemberRole">EventTypeArg.IsGroupChangeMemberRole</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsGroupChangeMemberRole">EventTypeArg.AsGroupChangeMemberRole</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsGroupCreate">EventTypeArg.IsGroupCreate</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsGroupCreate">EventTypeArg.AsGroupCreate</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsGroupDelete">EventTypeArg.IsGroupDelete</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsGroupDelete">EventTypeArg.AsGroupDelete</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsGroupDescriptionUpdated">EventTypeArg.IsGroupDescriptionUpdated</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsGroupDescriptionUpdated">EventTypeArg.AsGroupDescriptionUpdated</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsGroupJoinPolicyUpdated">EventTypeArg.IsGroupJoinPolicyUpdated</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsGroupJoinPolicyUpdated">EventTypeArg.AsGroupJoinPolicyUpdated</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsGroupMoved">EventTypeArg.IsGroupMoved</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsGroupMoved">EventTypeArg.AsGroupMoved</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsGroupRemoveExternalId">EventTypeArg.IsGroupRemoveExternalId</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsGroupRemoveExternalId">EventTypeArg.AsGroupRemoveExternalId</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsGroupRemoveMember">EventTypeArg.IsGroupRemoveMember</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsGroupRemoveMember">EventTypeArg.AsGroupRemoveMember</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsGroupRename">EventTypeArg.IsGroupRename</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsGroupRename">EventTypeArg.AsGroupRename</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsAccountLockOrUnlocked">EventTypeArg.IsAccountLockOrUnlocked</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsAccountLockOrUnlocked">EventTypeArg.AsAccountLockOrUnlocked</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsEmmError">EventTypeArg.IsEmmError</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsEmmError">EventTypeArg.AsEmmError</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsGuestAdminSignedInViaTrustedTeams">EventTypeArg.IsGuestAdminSignedInViaTrustedTeams</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsGuestAdminSignedInViaTrustedTeams">EventTypeArg.AsGuestAdminSignedInViaTrustedTeams</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsGuestAdminSignedOutViaTrustedTeams">EventTypeArg.IsGuestAdminSignedOutViaTrustedTeams</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsGuestAdminSignedOutViaTrustedTeams">EventTypeArg.AsGuestAdminSignedOutViaTrustedTeams</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsLoginFail">EventTypeArg.IsLoginFail</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsLoginFail">EventTypeArg.AsLoginFail</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsLoginSuccess">EventTypeArg.IsLoginSuccess</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsLoginSuccess">EventTypeArg.AsLoginSuccess</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsLogout">EventTypeArg.IsLogout</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsLogout">EventTypeArg.AsLogout</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsResellerSupportSessionEnd">EventTypeArg.IsResellerSupportSessionEnd</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsResellerSupportSessionEnd">EventTypeArg.AsResellerSupportSessionEnd</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsResellerSupportSessionStart">EventTypeArg.IsResellerSupportSessionStart</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsResellerSupportSessionStart">EventTypeArg.AsResellerSupportSessionStart</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSignInAsSessionEnd">EventTypeArg.IsSignInAsSessionEnd</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSignInAsSessionEnd">EventTypeArg.AsSignInAsSessionEnd</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSignInAsSessionStart">EventTypeArg.IsSignInAsSessionStart</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSignInAsSessionStart">EventTypeArg.AsSignInAsSessionStart</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSsoError">EventTypeArg.IsSsoError</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSsoError">EventTypeArg.AsSsoError</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsCreateTeamInviteLink">EventTypeArg.IsCreateTeamInviteLink</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsCreateTeamInviteLink">EventTypeArg.AsCreateTeamInviteLink</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDeleteTeamInviteLink">EventTypeArg.IsDeleteTeamInviteLink</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDeleteTeamInviteLink">EventTypeArg.AsDeleteTeamInviteLink</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsMemberAddExternalId">EventTypeArg.IsMemberAddExternalId</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsMemberAddExternalId">EventTypeArg.AsMemberAddExternalId</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsMemberAddName">EventTypeArg.IsMemberAddName</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsMemberAddName">EventTypeArg.AsMemberAddName</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsMemberChangeAdminRole">EventTypeArg.IsMemberChangeAdminRole</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsMemberChangeAdminRole">EventTypeArg.AsMemberChangeAdminRole</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsMemberChangeEmail">EventTypeArg.IsMemberChangeEmail</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsMemberChangeEmail">EventTypeArg.AsMemberChangeEmail</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsMemberChangeExternalId">EventTypeArg.IsMemberChangeExternalId</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsMemberChangeExternalId">EventTypeArg.AsMemberChangeExternalId</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsMemberChangeMembershipType">EventTypeArg.IsMemberChangeMembershipType</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsMemberChangeMembershipType">EventTypeArg.AsMemberChangeMembershipType</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsMemberChangeName">EventTypeArg.IsMemberChangeName</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsMemberChangeName">EventTypeArg.AsMemberChangeName</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsMemberChangeResellerRole">EventTypeArg.IsMemberChangeResellerRole</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsMemberChangeResellerRole">EventTypeArg.AsMemberChangeResellerRole</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsMemberChangeStatus">EventTypeArg.IsMemberChangeStatus</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsMemberChangeStatus">EventTypeArg.AsMemberChangeStatus</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsMemberDeleteManualContacts">EventTypeArg.IsMemberDeleteManualContacts</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsMemberDeleteManualContacts">EventTypeArg.AsMemberDeleteManualContacts</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsMemberDeleteProfilePhoto">EventTypeArg.IsMemberDeleteProfilePhoto</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsMemberDeleteProfilePhoto">EventTypeArg.AsMemberDeleteProfilePhoto</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsMemberPermanentlyDeleteAccountContents">EventTypeArg.IsMemberPermanentlyDeleteAccountContents</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsMemberPermanentlyDeleteAccountContents">EventTypeArg.AsMemberPermanentlyDeleteAccountContents</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsMemberRemoveExternalId">EventTypeArg.IsMemberRemoveExternalId</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsMemberRemoveExternalId">EventTypeArg.AsMemberRemoveExternalId</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsMemberSetProfilePhoto">EventTypeArg.IsMemberSetProfilePhoto</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsMemberSetProfilePhoto">EventTypeArg.AsMemberSetProfilePhoto</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsMemberSpaceLimitsAddCustomQuota">EventTypeArg.IsMemberSpaceLimitsAddCustomQuota</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsMemberSpaceLimitsAddCustomQuota">EventTypeArg.AsMemberSpaceLimitsAddCustomQuota</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsMemberSpaceLimitsChangeCustomQuota">EventTypeArg.IsMemberSpaceLimitsChangeCustomQuota</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsMemberSpaceLimitsChangeCustomQuota">EventTypeArg.AsMemberSpaceLimitsChangeCustomQuota</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsMemberSpaceLimitsChangeStatus">EventTypeArg.IsMemberSpaceLimitsChangeStatus</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsMemberSpaceLimitsChangeStatus">EventTypeArg.AsMemberSpaceLimitsChangeStatus</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsMemberSpaceLimitsRemoveCustomQuota">EventTypeArg.IsMemberSpaceLimitsRemoveCustomQuota</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsMemberSpaceLimitsRemoveCustomQuota">EventTypeArg.AsMemberSpaceLimitsRemoveCustomQuota</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsMemberSuggest">EventTypeArg.IsMemberSuggest</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsMemberSuggest">EventTypeArg.AsMemberSuggest</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsMemberTransferAccountContents">EventTypeArg.IsMemberTransferAccountContents</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsMemberTransferAccountContents">EventTypeArg.AsMemberTransferAccountContents</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPendingSecondaryEmailAdded">EventTypeArg.IsPendingSecondaryEmailAdded</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPendingSecondaryEmailAdded">EventTypeArg.AsPendingSecondaryEmailAdded</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSecondaryEmailDeleted">EventTypeArg.IsSecondaryEmailDeleted</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSecondaryEmailDeleted">EventTypeArg.AsSecondaryEmailDeleted</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSecondaryEmailVerified">EventTypeArg.IsSecondaryEmailVerified</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSecondaryEmailVerified">EventTypeArg.AsSecondaryEmailVerified</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSecondaryMailsPolicyChanged">EventTypeArg.IsSecondaryMailsPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSecondaryMailsPolicyChanged">EventTypeArg.AsSecondaryMailsPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsBinderAddPage">EventTypeArg.IsBinderAddPage</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsBinderAddPage">EventTypeArg.AsBinderAddPage</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsBinderAddSection">EventTypeArg.IsBinderAddSection</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsBinderAddSection">EventTypeArg.AsBinderAddSection</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsBinderRemovePage">EventTypeArg.IsBinderRemovePage</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsBinderRemovePage">EventTypeArg.AsBinderRemovePage</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsBinderRemoveSection">EventTypeArg.IsBinderRemoveSection</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsBinderRemoveSection">EventTypeArg.AsBinderRemoveSection</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsBinderRenamePage">EventTypeArg.IsBinderRenamePage</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsBinderRenamePage">EventTypeArg.AsBinderRenamePage</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsBinderRenameSection">EventTypeArg.IsBinderRenameSection</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsBinderRenameSection">EventTypeArg.AsBinderRenameSection</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsBinderReorderPage">EventTypeArg.IsBinderReorderPage</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsBinderReorderPage">EventTypeArg.AsBinderReorderPage</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsBinderReorderSection">EventTypeArg.IsBinderReorderSection</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsBinderReorderSection">EventTypeArg.AsBinderReorderSection</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperContentAddMember">EventTypeArg.IsPaperContentAddMember</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperContentAddMember">EventTypeArg.AsPaperContentAddMember</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperContentAddToFolder">EventTypeArg.IsPaperContentAddToFolder</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperContentAddToFolder">EventTypeArg.AsPaperContentAddToFolder</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperContentArchive">EventTypeArg.IsPaperContentArchive</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperContentArchive">EventTypeArg.AsPaperContentArchive</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperContentCreate">EventTypeArg.IsPaperContentCreate</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperContentCreate">EventTypeArg.AsPaperContentCreate</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperContentPermanentlyDelete">EventTypeArg.IsPaperContentPermanentlyDelete</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperContentPermanentlyDelete">EventTypeArg.AsPaperContentPermanentlyDelete</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperContentRemoveFromFolder">EventTypeArg.IsPaperContentRemoveFromFolder</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperContentRemoveFromFolder">EventTypeArg.AsPaperContentRemoveFromFolder</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperContentRemoveMember">EventTypeArg.IsPaperContentRemoveMember</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperContentRemoveMember">EventTypeArg.AsPaperContentRemoveMember</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperContentRename">EventTypeArg.IsPaperContentRename</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperContentRename">EventTypeArg.AsPaperContentRename</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperContentRestore">EventTypeArg.IsPaperContentRestore</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperContentRestore">EventTypeArg.AsPaperContentRestore</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperDocAddComment">EventTypeArg.IsPaperDocAddComment</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperDocAddComment">EventTypeArg.AsPaperDocAddComment</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperDocChangeMemberRole">EventTypeArg.IsPaperDocChangeMemberRole</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperDocChangeMemberRole">EventTypeArg.AsPaperDocChangeMemberRole</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperDocChangeSharingPolicy">EventTypeArg.IsPaperDocChangeSharingPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperDocChangeSharingPolicy">EventTypeArg.AsPaperDocChangeSharingPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperDocChangeSubscription">EventTypeArg.IsPaperDocChangeSubscription</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperDocChangeSubscription">EventTypeArg.AsPaperDocChangeSubscription</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperDocDeleted">EventTypeArg.IsPaperDocDeleted</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperDocDeleted">EventTypeArg.AsPaperDocDeleted</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperDocDeleteComment">EventTypeArg.IsPaperDocDeleteComment</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperDocDeleteComment">EventTypeArg.AsPaperDocDeleteComment</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperDocDownload">EventTypeArg.IsPaperDocDownload</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperDocDownload">EventTypeArg.AsPaperDocDownload</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperDocEdit">EventTypeArg.IsPaperDocEdit</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperDocEdit">EventTypeArg.AsPaperDocEdit</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperDocEditComment">EventTypeArg.IsPaperDocEditComment</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperDocEditComment">EventTypeArg.AsPaperDocEditComment</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperDocFollowed">EventTypeArg.IsPaperDocFollowed</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperDocFollowed">EventTypeArg.AsPaperDocFollowed</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperDocMention">EventTypeArg.IsPaperDocMention</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperDocMention">EventTypeArg.AsPaperDocMention</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperDocOwnershipChanged">EventTypeArg.IsPaperDocOwnershipChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperDocOwnershipChanged">EventTypeArg.AsPaperDocOwnershipChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperDocRequestAccess">EventTypeArg.IsPaperDocRequestAccess</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperDocRequestAccess">EventTypeArg.AsPaperDocRequestAccess</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperDocResolveComment">EventTypeArg.IsPaperDocResolveComment</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperDocResolveComment">EventTypeArg.AsPaperDocResolveComment</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperDocRevert">EventTypeArg.IsPaperDocRevert</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperDocRevert">EventTypeArg.AsPaperDocRevert</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperDocSlackShare">EventTypeArg.IsPaperDocSlackShare</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperDocSlackShare">EventTypeArg.AsPaperDocSlackShare</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperDocTeamInvite">EventTypeArg.IsPaperDocTeamInvite</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperDocTeamInvite">EventTypeArg.AsPaperDocTeamInvite</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperDocTrashed">EventTypeArg.IsPaperDocTrashed</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperDocTrashed">EventTypeArg.AsPaperDocTrashed</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperDocUnresolveComment">EventTypeArg.IsPaperDocUnresolveComment</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperDocUnresolveComment">EventTypeArg.AsPaperDocUnresolveComment</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperDocUntrashed">EventTypeArg.IsPaperDocUntrashed</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperDocUntrashed">EventTypeArg.AsPaperDocUntrashed</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperDocView">EventTypeArg.IsPaperDocView</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperDocView">EventTypeArg.AsPaperDocView</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperExternalViewAllow">EventTypeArg.IsPaperExternalViewAllow</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperExternalViewAllow">EventTypeArg.AsPaperExternalViewAllow</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperExternalViewDefaultTeam">EventTypeArg.IsPaperExternalViewDefaultTeam</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperExternalViewDefaultTeam">EventTypeArg.AsPaperExternalViewDefaultTeam</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperExternalViewForbid">EventTypeArg.IsPaperExternalViewForbid</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperExternalViewForbid">EventTypeArg.AsPaperExternalViewForbid</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperFolderChangeSubscription">EventTypeArg.IsPaperFolderChangeSubscription</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperFolderChangeSubscription">EventTypeArg.AsPaperFolderChangeSubscription</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperFolderDeleted">EventTypeArg.IsPaperFolderDeleted</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperFolderDeleted">EventTypeArg.AsPaperFolderDeleted</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperFolderFollowed">EventTypeArg.IsPaperFolderFollowed</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperFolderFollowed">EventTypeArg.AsPaperFolderFollowed</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperFolderTeamInvite">EventTypeArg.IsPaperFolderTeamInvite</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperFolderTeamInvite">EventTypeArg.AsPaperFolderTeamInvite</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperPublishedLinkChangePermission">EventTypeArg.IsPaperPublishedLinkChangePermission</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperPublishedLinkChangePermission">EventTypeArg.AsPaperPublishedLinkChangePermission</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperPublishedLinkCreate">EventTypeArg.IsPaperPublishedLinkCreate</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperPublishedLinkCreate">EventTypeArg.AsPaperPublishedLinkCreate</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperPublishedLinkDisabled">EventTypeArg.IsPaperPublishedLinkDisabled</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperPublishedLinkDisabled">EventTypeArg.AsPaperPublishedLinkDisabled</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperPublishedLinkView">EventTypeArg.IsPaperPublishedLinkView</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperPublishedLinkView">EventTypeArg.AsPaperPublishedLinkView</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPasswordChange">EventTypeArg.IsPasswordChange</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPasswordChange">EventTypeArg.AsPasswordChange</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPasswordReset">EventTypeArg.IsPasswordReset</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPasswordReset">EventTypeArg.AsPasswordReset</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPasswordResetAll">EventTypeArg.IsPasswordResetAll</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPasswordResetAll">EventTypeArg.AsPasswordResetAll</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsClassificationCreateReport">EventTypeArg.IsClassificationCreateReport</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsClassificationCreateReport">EventTypeArg.AsClassificationCreateReport</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsClassificationCreateReportFail">EventTypeArg.IsClassificationCreateReportFail</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsClassificationCreateReportFail">EventTypeArg.AsClassificationCreateReportFail</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsEmmCreateExceptionsReport">EventTypeArg.IsEmmCreateExceptionsReport</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsEmmCreateExceptionsReport">EventTypeArg.AsEmmCreateExceptionsReport</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsEmmCreateUsageReport">EventTypeArg.IsEmmCreateUsageReport</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsEmmCreateUsageReport">EventTypeArg.AsEmmCreateUsageReport</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsExportMembersReport">EventTypeArg.IsExportMembersReport</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsExportMembersReport">EventTypeArg.AsExportMembersReport</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsExportMembersReportFail">EventTypeArg.IsExportMembersReportFail</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsExportMembersReportFail">EventTypeArg.AsExportMembersReportFail</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsExternalSharingCreateReport">EventTypeArg.IsExternalSharingCreateReport</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsExternalSharingCreateReport">EventTypeArg.AsExternalSharingCreateReport</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsExternalSharingReportFailed">EventTypeArg.IsExternalSharingReportFailed</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsExternalSharingReportFailed">EventTypeArg.AsExternalSharingReportFailed</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsNoExpirationLinkGenCreateReport">EventTypeArg.IsNoExpirationLinkGenCreateReport</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsNoExpirationLinkGenCreateReport">EventTypeArg.AsNoExpirationLinkGenCreateReport</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsNoExpirationLinkGenReportFailed">EventTypeArg.IsNoExpirationLinkGenReportFailed</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsNoExpirationLinkGenReportFailed">EventTypeArg.AsNoExpirationLinkGenReportFailed</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsNoPasswordLinkGenCreateReport">EventTypeArg.IsNoPasswordLinkGenCreateReport</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsNoPasswordLinkGenCreateReport">EventTypeArg.AsNoPasswordLinkGenCreateReport</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsNoPasswordLinkGenReportFailed">EventTypeArg.IsNoPasswordLinkGenReportFailed</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsNoPasswordLinkGenReportFailed">EventTypeArg.AsNoPasswordLinkGenReportFailed</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsNoPasswordLinkViewCreateReport">EventTypeArg.IsNoPasswordLinkViewCreateReport</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsNoPasswordLinkViewCreateReport">EventTypeArg.AsNoPasswordLinkViewCreateReport</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsNoPasswordLinkViewReportFailed">EventTypeArg.IsNoPasswordLinkViewReportFailed</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsNoPasswordLinkViewReportFailed">EventTypeArg.AsNoPasswordLinkViewReportFailed</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsOutdatedLinkViewCreateReport">EventTypeArg.IsOutdatedLinkViewCreateReport</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsOutdatedLinkViewCreateReport">EventTypeArg.AsOutdatedLinkViewCreateReport</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsOutdatedLinkViewReportFailed">EventTypeArg.IsOutdatedLinkViewReportFailed</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsOutdatedLinkViewReportFailed">EventTypeArg.AsOutdatedLinkViewReportFailed</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperAdminExportStart">EventTypeArg.IsPaperAdminExportStart</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperAdminExportStart">EventTypeArg.AsPaperAdminExportStart</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSmartSyncCreateAdminPrivilegeReport">EventTypeArg.IsSmartSyncCreateAdminPrivilegeReport</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSmartSyncCreateAdminPrivilegeReport">EventTypeArg.AsSmartSyncCreateAdminPrivilegeReport</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamActivityCreateReport">EventTypeArg.IsTeamActivityCreateReport</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamActivityCreateReport">EventTypeArg.AsTeamActivityCreateReport</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamActivityCreateReportFail">EventTypeArg.IsTeamActivityCreateReportFail</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamActivityCreateReportFail">EventTypeArg.AsTeamActivityCreateReportFail</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsCollectionShare">EventTypeArg.IsCollectionShare</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsCollectionShare">EventTypeArg.AsCollectionShare</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileTransfersFileAdd">EventTypeArg.IsFileTransfersFileAdd</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileTransfersFileAdd">EventTypeArg.AsFileTransfersFileAdd</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileTransfersTransferDelete">EventTypeArg.IsFileTransfersTransferDelete</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileTransfersTransferDelete">EventTypeArg.AsFileTransfersTransferDelete</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileTransfersTransferDownload">EventTypeArg.IsFileTransfersTransferDownload</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileTransfersTransferDownload">EventTypeArg.AsFileTransfersTransferDownload</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileTransfersTransferSend">EventTypeArg.IsFileTransfersTransferSend</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileTransfersTransferSend">EventTypeArg.AsFileTransfersTransferSend</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileTransfersTransferView">EventTypeArg.IsFileTransfersTransferView</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileTransfersTransferView">EventTypeArg.AsFileTransfersTransferView</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsNoteAclInviteOnly">EventTypeArg.IsNoteAclInviteOnly</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsNoteAclInviteOnly">EventTypeArg.AsNoteAclInviteOnly</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsNoteAclLink">EventTypeArg.IsNoteAclLink</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsNoteAclLink">EventTypeArg.AsNoteAclLink</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsNoteAclTeamLink">EventTypeArg.IsNoteAclTeamLink</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsNoteAclTeamLink">EventTypeArg.AsNoteAclTeamLink</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsNoteShared">EventTypeArg.IsNoteShared</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsNoteShared">EventTypeArg.AsNoteShared</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsNoteShareReceive">EventTypeArg.IsNoteShareReceive</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsNoteShareReceive">EventTypeArg.AsNoteShareReceive</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsOpenNoteShared">EventTypeArg.IsOpenNoteShared</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsOpenNoteShared">EventTypeArg.AsOpenNoteShared</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSfAddGroup">EventTypeArg.IsSfAddGroup</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSfAddGroup">EventTypeArg.AsSfAddGroup</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSfAllowNonMembersToViewSharedLinks">EventTypeArg.IsSfAllowNonMembersToViewSharedLinks</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSfAllowNonMembersToViewSharedLinks">EventTypeArg.AsSfAllowNonMembersToViewSharedLinks</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSfExternalInviteWarn">EventTypeArg.IsSfExternalInviteWarn</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSfExternalInviteWarn">EventTypeArg.AsSfExternalInviteWarn</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSfFbInvite">EventTypeArg.IsSfFbInvite</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSfFbInvite">EventTypeArg.AsSfFbInvite</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSfFbInviteChangeRole">EventTypeArg.IsSfFbInviteChangeRole</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSfFbInviteChangeRole">EventTypeArg.AsSfFbInviteChangeRole</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSfFbUninvite">EventTypeArg.IsSfFbUninvite</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSfFbUninvite">EventTypeArg.AsSfFbUninvite</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSfInviteGroup">EventTypeArg.IsSfInviteGroup</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSfInviteGroup">EventTypeArg.AsSfInviteGroup</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSfTeamGrantAccess">EventTypeArg.IsSfTeamGrantAccess</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSfTeamGrantAccess">EventTypeArg.AsSfTeamGrantAccess</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSfTeamInvite">EventTypeArg.IsSfTeamInvite</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSfTeamInvite">EventTypeArg.AsSfTeamInvite</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSfTeamInviteChangeRole">EventTypeArg.IsSfTeamInviteChangeRole</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSfTeamInviteChangeRole">EventTypeArg.AsSfTeamInviteChangeRole</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSfTeamJoin">EventTypeArg.IsSfTeamJoin</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSfTeamJoin">EventTypeArg.AsSfTeamJoin</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSfTeamJoinFromOobLink">EventTypeArg.IsSfTeamJoinFromOobLink</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSfTeamJoinFromOobLink">EventTypeArg.AsSfTeamJoinFromOobLink</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSfTeamUninvite">EventTypeArg.IsSfTeamUninvite</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSfTeamUninvite">EventTypeArg.AsSfTeamUninvite</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedContentAddInvitees">EventTypeArg.IsSharedContentAddInvitees</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedContentAddInvitees">EventTypeArg.AsSharedContentAddInvitees</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedContentAddLinkExpiry">EventTypeArg.IsSharedContentAddLinkExpiry</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedContentAddLinkExpiry">EventTypeArg.AsSharedContentAddLinkExpiry</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedContentAddLinkPassword">EventTypeArg.IsSharedContentAddLinkPassword</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedContentAddLinkPassword">EventTypeArg.AsSharedContentAddLinkPassword</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedContentAddMember">EventTypeArg.IsSharedContentAddMember</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedContentAddMember">EventTypeArg.AsSharedContentAddMember</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedContentChangeDownloadsPolicy">EventTypeArg.IsSharedContentChangeDownloadsPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedContentChangeDownloadsPolicy">EventTypeArg.AsSharedContentChangeDownloadsPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedContentChangeInviteeRole">EventTypeArg.IsSharedContentChangeInviteeRole</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedContentChangeInviteeRole">EventTypeArg.AsSharedContentChangeInviteeRole</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedContentChangeLinkAudience">EventTypeArg.IsSharedContentChangeLinkAudience</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedContentChangeLinkAudience">EventTypeArg.AsSharedContentChangeLinkAudience</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedContentChangeLinkExpiry">EventTypeArg.IsSharedContentChangeLinkExpiry</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedContentChangeLinkExpiry">EventTypeArg.AsSharedContentChangeLinkExpiry</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedContentChangeLinkPassword">EventTypeArg.IsSharedContentChangeLinkPassword</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedContentChangeLinkPassword">EventTypeArg.AsSharedContentChangeLinkPassword</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedContentChangeMemberRole">EventTypeArg.IsSharedContentChangeMemberRole</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedContentChangeMemberRole">EventTypeArg.AsSharedContentChangeMemberRole</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedContentChangeViewerInfoPolicy">EventTypeArg.IsSharedContentChangeViewerInfoPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedContentChangeViewerInfoPolicy">EventTypeArg.AsSharedContentChangeViewerInfoPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedContentClaimInvitation">EventTypeArg.IsSharedContentClaimInvitation</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedContentClaimInvitation">EventTypeArg.AsSharedContentClaimInvitation</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedContentCopy">EventTypeArg.IsSharedContentCopy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedContentCopy">EventTypeArg.AsSharedContentCopy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedContentDownload">EventTypeArg.IsSharedContentDownload</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedContentDownload">EventTypeArg.AsSharedContentDownload</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedContentRelinquishMembership">EventTypeArg.IsSharedContentRelinquishMembership</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedContentRelinquishMembership">EventTypeArg.AsSharedContentRelinquishMembership</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedContentRemoveInvitees">EventTypeArg.IsSharedContentRemoveInvitees</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedContentRemoveInvitees">EventTypeArg.AsSharedContentRemoveInvitees</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedContentRemoveLinkExpiry">EventTypeArg.IsSharedContentRemoveLinkExpiry</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedContentRemoveLinkExpiry">EventTypeArg.AsSharedContentRemoveLinkExpiry</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedContentRemoveLinkPassword">EventTypeArg.IsSharedContentRemoveLinkPassword</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedContentRemoveLinkPassword">EventTypeArg.AsSharedContentRemoveLinkPassword</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedContentRemoveMember">EventTypeArg.IsSharedContentRemoveMember</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedContentRemoveMember">EventTypeArg.AsSharedContentRemoveMember</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedContentRequestAccess">EventTypeArg.IsSharedContentRequestAccess</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedContentRequestAccess">EventTypeArg.AsSharedContentRequestAccess</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedContentRestoreInvitees">EventTypeArg.IsSharedContentRestoreInvitees</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedContentRestoreInvitees">EventTypeArg.AsSharedContentRestoreInvitees</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedContentRestoreMember">EventTypeArg.IsSharedContentRestoreMember</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedContentRestoreMember">EventTypeArg.AsSharedContentRestoreMember</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedContentUnshare">EventTypeArg.IsSharedContentUnshare</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedContentUnshare">EventTypeArg.AsSharedContentUnshare</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedContentView">EventTypeArg.IsSharedContentView</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedContentView">EventTypeArg.AsSharedContentView</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedFolderChangeLinkPolicy">EventTypeArg.IsSharedFolderChangeLinkPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedFolderChangeLinkPolicy">EventTypeArg.AsSharedFolderChangeLinkPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedFolderChangeMembersInheritancePolicy">EventTypeArg.IsSharedFolderChangeMembersInheritancePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedFolderChangeMembersInheritancePolicy">EventTypeArg.AsSharedFolderChangeMembersInheritancePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedFolderChangeMembersManagementPolicy">EventTypeArg.IsSharedFolderChangeMembersManagementPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedFolderChangeMembersManagementPolicy">EventTypeArg.AsSharedFolderChangeMembersManagementPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedFolderChangeMembersPolicy">EventTypeArg.IsSharedFolderChangeMembersPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedFolderChangeMembersPolicy">EventTypeArg.AsSharedFolderChangeMembersPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedFolderCreate">EventTypeArg.IsSharedFolderCreate</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedFolderCreate">EventTypeArg.AsSharedFolderCreate</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedFolderDeclineInvitation">EventTypeArg.IsSharedFolderDeclineInvitation</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedFolderDeclineInvitation">EventTypeArg.AsSharedFolderDeclineInvitation</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedFolderMount">EventTypeArg.IsSharedFolderMount</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedFolderMount">EventTypeArg.AsSharedFolderMount</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedFolderNest">EventTypeArg.IsSharedFolderNest</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedFolderNest">EventTypeArg.AsSharedFolderNest</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedFolderTransferOwnership">EventTypeArg.IsSharedFolderTransferOwnership</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedFolderTransferOwnership">EventTypeArg.AsSharedFolderTransferOwnership</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedFolderUnmount">EventTypeArg.IsSharedFolderUnmount</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedFolderUnmount">EventTypeArg.AsSharedFolderUnmount</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedLinkAddExpiry">EventTypeArg.IsSharedLinkAddExpiry</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedLinkAddExpiry">EventTypeArg.AsSharedLinkAddExpiry</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedLinkChangeExpiry">EventTypeArg.IsSharedLinkChangeExpiry</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedLinkChangeExpiry">EventTypeArg.AsSharedLinkChangeExpiry</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedLinkChangeVisibility">EventTypeArg.IsSharedLinkChangeVisibility</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedLinkChangeVisibility">EventTypeArg.AsSharedLinkChangeVisibility</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedLinkCopy">EventTypeArg.IsSharedLinkCopy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedLinkCopy">EventTypeArg.AsSharedLinkCopy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedLinkCreate">EventTypeArg.IsSharedLinkCreate</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedLinkCreate">EventTypeArg.AsSharedLinkCreate</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedLinkDisable">EventTypeArg.IsSharedLinkDisable</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedLinkDisable">EventTypeArg.AsSharedLinkDisable</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedLinkDownload">EventTypeArg.IsSharedLinkDownload</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedLinkDownload">EventTypeArg.AsSharedLinkDownload</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedLinkRemoveExpiry">EventTypeArg.IsSharedLinkRemoveExpiry</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedLinkRemoveExpiry">EventTypeArg.AsSharedLinkRemoveExpiry</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedLinkSettingsAddExpiration">EventTypeArg.IsSharedLinkSettingsAddExpiration</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedLinkSettingsAddExpiration">EventTypeArg.AsSharedLinkSettingsAddExpiration</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedLinkSettingsAddPassword">EventTypeArg.IsSharedLinkSettingsAddPassword</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedLinkSettingsAddPassword">EventTypeArg.AsSharedLinkSettingsAddPassword</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedLinkSettingsAllowDownloadDisabled">EventTypeArg.IsSharedLinkSettingsAllowDownloadDisabled</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedLinkSettingsAllowDownloadDisabled">EventTypeArg.AsSharedLinkSettingsAllowDownloadDisabled</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedLinkSettingsAllowDownloadEnabled">EventTypeArg.IsSharedLinkSettingsAllowDownloadEnabled</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedLinkSettingsAllowDownloadEnabled">EventTypeArg.AsSharedLinkSettingsAllowDownloadEnabled</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedLinkSettingsChangeAudience">EventTypeArg.IsSharedLinkSettingsChangeAudience</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedLinkSettingsChangeAudience">EventTypeArg.AsSharedLinkSettingsChangeAudience</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedLinkSettingsChangeExpiration">EventTypeArg.IsSharedLinkSettingsChangeExpiration</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedLinkSettingsChangeExpiration">EventTypeArg.AsSharedLinkSettingsChangeExpiration</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedLinkSettingsChangePassword">EventTypeArg.IsSharedLinkSettingsChangePassword</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedLinkSettingsChangePassword">EventTypeArg.AsSharedLinkSettingsChangePassword</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedLinkSettingsRemoveExpiration">EventTypeArg.IsSharedLinkSettingsRemoveExpiration</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedLinkSettingsRemoveExpiration">EventTypeArg.AsSharedLinkSettingsRemoveExpiration</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedLinkSettingsRemovePassword">EventTypeArg.IsSharedLinkSettingsRemovePassword</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedLinkSettingsRemovePassword">EventTypeArg.AsSharedLinkSettingsRemovePassword</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedLinkShare">EventTypeArg.IsSharedLinkShare</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedLinkShare">EventTypeArg.AsSharedLinkShare</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedLinkView">EventTypeArg.IsSharedLinkView</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedLinkView">EventTypeArg.AsSharedLinkView</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharedNoteOpened">EventTypeArg.IsSharedNoteOpened</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharedNoteOpened">EventTypeArg.AsSharedNoteOpened</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsShmodelDisableDownloads">EventTypeArg.IsShmodelDisableDownloads</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsShmodelDisableDownloads">EventTypeArg.AsShmodelDisableDownloads</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsShmodelEnableDownloads">EventTypeArg.IsShmodelEnableDownloads</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsShmodelEnableDownloads">EventTypeArg.AsShmodelEnableDownloads</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsShmodelGroupShare">EventTypeArg.IsShmodelGroupShare</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsShmodelGroupShare">EventTypeArg.AsShmodelGroupShare</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsShowcaseAccessGranted">EventTypeArg.IsShowcaseAccessGranted</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsShowcaseAccessGranted">EventTypeArg.AsShowcaseAccessGranted</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsShowcaseAddMember">EventTypeArg.IsShowcaseAddMember</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsShowcaseAddMember">EventTypeArg.AsShowcaseAddMember</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsShowcaseArchived">EventTypeArg.IsShowcaseArchived</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsShowcaseArchived">EventTypeArg.AsShowcaseArchived</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsShowcaseCreated">EventTypeArg.IsShowcaseCreated</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsShowcaseCreated">EventTypeArg.AsShowcaseCreated</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsShowcaseDeleteComment">EventTypeArg.IsShowcaseDeleteComment</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsShowcaseDeleteComment">EventTypeArg.AsShowcaseDeleteComment</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsShowcaseEdited">EventTypeArg.IsShowcaseEdited</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsShowcaseEdited">EventTypeArg.AsShowcaseEdited</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsShowcaseEditComment">EventTypeArg.IsShowcaseEditComment</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsShowcaseEditComment">EventTypeArg.AsShowcaseEditComment</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsShowcaseFileAdded">EventTypeArg.IsShowcaseFileAdded</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsShowcaseFileAdded">EventTypeArg.AsShowcaseFileAdded</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsShowcaseFileDownload">EventTypeArg.IsShowcaseFileDownload</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsShowcaseFileDownload">EventTypeArg.AsShowcaseFileDownload</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsShowcaseFileRemoved">EventTypeArg.IsShowcaseFileRemoved</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsShowcaseFileRemoved">EventTypeArg.AsShowcaseFileRemoved</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsShowcaseFileView">EventTypeArg.IsShowcaseFileView</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsShowcaseFileView">EventTypeArg.AsShowcaseFileView</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsShowcasePermanentlyDeleted">EventTypeArg.IsShowcasePermanentlyDeleted</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsShowcasePermanentlyDeleted">EventTypeArg.AsShowcasePermanentlyDeleted</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsShowcasePostComment">EventTypeArg.IsShowcasePostComment</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsShowcasePostComment">EventTypeArg.AsShowcasePostComment</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsShowcaseRemoveMember">EventTypeArg.IsShowcaseRemoveMember</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsShowcaseRemoveMember">EventTypeArg.AsShowcaseRemoveMember</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsShowcaseRenamed">EventTypeArg.IsShowcaseRenamed</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsShowcaseRenamed">EventTypeArg.AsShowcaseRenamed</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsShowcaseRequestAccess">EventTypeArg.IsShowcaseRequestAccess</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsShowcaseRequestAccess">EventTypeArg.AsShowcaseRequestAccess</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsShowcaseResolveComment">EventTypeArg.IsShowcaseResolveComment</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsShowcaseResolveComment">EventTypeArg.AsShowcaseResolveComment</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsShowcaseRestored">EventTypeArg.IsShowcaseRestored</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsShowcaseRestored">EventTypeArg.AsShowcaseRestored</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsShowcaseTrashed">EventTypeArg.IsShowcaseTrashed</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsShowcaseTrashed">EventTypeArg.AsShowcaseTrashed</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsShowcaseTrashedDeprecated">EventTypeArg.IsShowcaseTrashedDeprecated</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsShowcaseTrashedDeprecated">EventTypeArg.AsShowcaseTrashedDeprecated</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsShowcaseUnresolveComment">EventTypeArg.IsShowcaseUnresolveComment</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsShowcaseUnresolveComment">EventTypeArg.AsShowcaseUnresolveComment</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsShowcaseUntrashed">EventTypeArg.IsShowcaseUntrashed</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsShowcaseUntrashed">EventTypeArg.AsShowcaseUntrashed</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsShowcaseUntrashedDeprecated">EventTypeArg.IsShowcaseUntrashedDeprecated</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsShowcaseUntrashedDeprecated">EventTypeArg.AsShowcaseUntrashedDeprecated</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsShowcaseView">EventTypeArg.IsShowcaseView</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsShowcaseView">EventTypeArg.AsShowcaseView</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSsoAddCert">EventTypeArg.IsSsoAddCert</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSsoAddCert">EventTypeArg.AsSsoAddCert</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSsoAddLoginUrl">EventTypeArg.IsSsoAddLoginUrl</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSsoAddLoginUrl">EventTypeArg.AsSsoAddLoginUrl</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSsoAddLogoutUrl">EventTypeArg.IsSsoAddLogoutUrl</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSsoAddLogoutUrl">EventTypeArg.AsSsoAddLogoutUrl</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSsoChangeCert">EventTypeArg.IsSsoChangeCert</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSsoChangeCert">EventTypeArg.AsSsoChangeCert</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSsoChangeLoginUrl">EventTypeArg.IsSsoChangeLoginUrl</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSsoChangeLoginUrl">EventTypeArg.AsSsoChangeLoginUrl</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSsoChangeLogoutUrl">EventTypeArg.IsSsoChangeLogoutUrl</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSsoChangeLogoutUrl">EventTypeArg.AsSsoChangeLogoutUrl</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSsoChangeSamlIdentityMode">EventTypeArg.IsSsoChangeSamlIdentityMode</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSsoChangeSamlIdentityMode">EventTypeArg.AsSsoChangeSamlIdentityMode</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSsoRemoveCert">EventTypeArg.IsSsoRemoveCert</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSsoRemoveCert">EventTypeArg.AsSsoRemoveCert</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSsoRemoveLoginUrl">EventTypeArg.IsSsoRemoveLoginUrl</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSsoRemoveLoginUrl">EventTypeArg.AsSsoRemoveLoginUrl</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSsoRemoveLogoutUrl">EventTypeArg.IsSsoRemoveLogoutUrl</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSsoRemoveLogoutUrl">EventTypeArg.AsSsoRemoveLogoutUrl</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamFolderChangeStatus">EventTypeArg.IsTeamFolderChangeStatus</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamFolderChangeStatus">EventTypeArg.AsTeamFolderChangeStatus</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamFolderCreate">EventTypeArg.IsTeamFolderCreate</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamFolderCreate">EventTypeArg.AsTeamFolderCreate</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamFolderDowngrade">EventTypeArg.IsTeamFolderDowngrade</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamFolderDowngrade">EventTypeArg.AsTeamFolderDowngrade</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamFolderPermanentlyDelete">EventTypeArg.IsTeamFolderPermanentlyDelete</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamFolderPermanentlyDelete">EventTypeArg.AsTeamFolderPermanentlyDelete</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamFolderRename">EventTypeArg.IsTeamFolderRename</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamFolderRename">EventTypeArg.AsTeamFolderRename</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamSelectiveSyncSettingsChanged">EventTypeArg.IsTeamSelectiveSyncSettingsChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamSelectiveSyncSettingsChanged">EventTypeArg.AsTeamSelectiveSyncSettingsChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsAccountCaptureChangePolicy">EventTypeArg.IsAccountCaptureChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsAccountCaptureChangePolicy">EventTypeArg.AsAccountCaptureChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsAllowDownloadDisabled">EventTypeArg.IsAllowDownloadDisabled</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsAllowDownloadDisabled">EventTypeArg.AsAllowDownloadDisabled</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsAllowDownloadEnabled">EventTypeArg.IsAllowDownloadEnabled</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsAllowDownloadEnabled">EventTypeArg.AsAllowDownloadEnabled</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsAppPermissionsChanged">EventTypeArg.IsAppPermissionsChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsAppPermissionsChanged">EventTypeArg.AsAppPermissionsChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsCameraUploadsPolicyChanged">EventTypeArg.IsCameraUploadsPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsCameraUploadsPolicyChanged">EventTypeArg.AsCameraUploadsPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsCaptureTranscriptPolicyChanged">EventTypeArg.IsCaptureTranscriptPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsCaptureTranscriptPolicyChanged">EventTypeArg.AsCaptureTranscriptPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsClassificationChangePolicy">EventTypeArg.IsClassificationChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsClassificationChangePolicy">EventTypeArg.AsClassificationChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsComputerBackupPolicyChanged">EventTypeArg.IsComputerBackupPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsComputerBackupPolicyChanged">EventTypeArg.AsComputerBackupPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsContentAdministrationPolicyChanged">EventTypeArg.IsContentAdministrationPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsContentAdministrationPolicyChanged">EventTypeArg.AsContentAdministrationPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDataPlacementRestrictionChangePolicy">EventTypeArg.IsDataPlacementRestrictionChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDataPlacementRestrictionChangePolicy">EventTypeArg.AsDataPlacementRestrictionChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDataPlacementRestrictionSatisfyPolicy">EventTypeArg.IsDataPlacementRestrictionSatisfyPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDataPlacementRestrictionSatisfyPolicy">EventTypeArg.AsDataPlacementRestrictionSatisfyPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDeviceApprovalsAddException">EventTypeArg.IsDeviceApprovalsAddException</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDeviceApprovalsAddException">EventTypeArg.AsDeviceApprovalsAddException</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDeviceApprovalsChangeDesktopPolicy">EventTypeArg.IsDeviceApprovalsChangeDesktopPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDeviceApprovalsChangeDesktopPolicy">EventTypeArg.AsDeviceApprovalsChangeDesktopPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDeviceApprovalsChangeMobilePolicy">EventTypeArg.IsDeviceApprovalsChangeMobilePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDeviceApprovalsChangeMobilePolicy">EventTypeArg.AsDeviceApprovalsChangeMobilePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDeviceApprovalsChangeOverageAction">EventTypeArg.IsDeviceApprovalsChangeOverageAction</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDeviceApprovalsChangeOverageAction">EventTypeArg.AsDeviceApprovalsChangeOverageAction</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDeviceApprovalsChangeUnlinkAction">EventTypeArg.IsDeviceApprovalsChangeUnlinkAction</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDeviceApprovalsChangeUnlinkAction">EventTypeArg.AsDeviceApprovalsChangeUnlinkAction</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDeviceApprovalsRemoveException">EventTypeArg.IsDeviceApprovalsRemoveException</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDeviceApprovalsRemoveException">EventTypeArg.AsDeviceApprovalsRemoveException</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDirectoryRestrictionsAddMembers">EventTypeArg.IsDirectoryRestrictionsAddMembers</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDirectoryRestrictionsAddMembers">EventTypeArg.AsDirectoryRestrictionsAddMembers</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDirectoryRestrictionsRemoveMembers">EventTypeArg.IsDirectoryRestrictionsRemoveMembers</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDirectoryRestrictionsRemoveMembers">EventTypeArg.AsDirectoryRestrictionsRemoveMembers</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDropboxPasswordsPolicyChanged">EventTypeArg.IsDropboxPasswordsPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDropboxPasswordsPolicyChanged">EventTypeArg.AsDropboxPasswordsPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsEmailIngestPolicyChanged">EventTypeArg.IsEmailIngestPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsEmailIngestPolicyChanged">EventTypeArg.AsEmailIngestPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsEmmAddException">EventTypeArg.IsEmmAddException</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsEmmAddException">EventTypeArg.AsEmmAddException</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsEmmChangePolicy">EventTypeArg.IsEmmChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsEmmChangePolicy">EventTypeArg.AsEmmChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsEmmRemoveException">EventTypeArg.IsEmmRemoveException</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsEmmRemoveException">EventTypeArg.AsEmmRemoveException</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsExtendedVersionHistoryChangePolicy">EventTypeArg.IsExtendedVersionHistoryChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsExtendedVersionHistoryChangePolicy">EventTypeArg.AsExtendedVersionHistoryChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsExternalDriveBackupPolicyChanged">EventTypeArg.IsExternalDriveBackupPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsExternalDriveBackupPolicyChanged">EventTypeArg.AsExternalDriveBackupPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileCommentsChangePolicy">EventTypeArg.IsFileCommentsChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileCommentsChangePolicy">EventTypeArg.AsFileCommentsChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileLockingPolicyChanged">EventTypeArg.IsFileLockingPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileLockingPolicyChanged">EventTypeArg.AsFileLockingPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileRequestsChangePolicy">EventTypeArg.IsFileRequestsChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileRequestsChangePolicy">EventTypeArg.AsFileRequestsChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileRequestsEmailsEnabled">EventTypeArg.IsFileRequestsEmailsEnabled</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileRequestsEmailsEnabled">EventTypeArg.AsFileRequestsEmailsEnabled</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileRequestsEmailsRestrictedToTeamOnly">EventTypeArg.IsFileRequestsEmailsRestrictedToTeamOnly</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileRequestsEmailsRestrictedToTeamOnly">EventTypeArg.AsFileRequestsEmailsRestrictedToTeamOnly</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsFileTransfersPolicyChanged">EventTypeArg.IsFileTransfersPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsFileTransfersPolicyChanged">EventTypeArg.AsFileTransfersPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsGoogleSsoChangePolicy">EventTypeArg.IsGoogleSsoChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsGoogleSsoChangePolicy">EventTypeArg.AsGoogleSsoChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsGroupUserManagementChangePolicy">EventTypeArg.IsGroupUserManagementChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsGroupUserManagementChangePolicy">EventTypeArg.AsGroupUserManagementChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsIntegrationPolicyChanged">EventTypeArg.IsIntegrationPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsIntegrationPolicyChanged">EventTypeArg.AsIntegrationPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsInviteAcceptanceEmailPolicyChanged">EventTypeArg.IsInviteAcceptanceEmailPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsInviteAcceptanceEmailPolicyChanged">EventTypeArg.AsInviteAcceptanceEmailPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsMemberRequestsChangePolicy">EventTypeArg.IsMemberRequestsChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsMemberRequestsChangePolicy">EventTypeArg.AsMemberRequestsChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsMemberSendInvitePolicyChanged">EventTypeArg.IsMemberSendInvitePolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsMemberSendInvitePolicyChanged">EventTypeArg.AsMemberSendInvitePolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsMemberSpaceLimitsAddException">EventTypeArg.IsMemberSpaceLimitsAddException</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsMemberSpaceLimitsAddException">EventTypeArg.AsMemberSpaceLimitsAddException</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsMemberSpaceLimitsChangeCapsTypePolicy">EventTypeArg.IsMemberSpaceLimitsChangeCapsTypePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsMemberSpaceLimitsChangeCapsTypePolicy">EventTypeArg.AsMemberSpaceLimitsChangeCapsTypePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsMemberSpaceLimitsChangePolicy">EventTypeArg.IsMemberSpaceLimitsChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsMemberSpaceLimitsChangePolicy">EventTypeArg.AsMemberSpaceLimitsChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsMemberSpaceLimitsRemoveException">EventTypeArg.IsMemberSpaceLimitsRemoveException</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsMemberSpaceLimitsRemoveException">EventTypeArg.AsMemberSpaceLimitsRemoveException</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsMemberSuggestionsChangePolicy">EventTypeArg.IsMemberSuggestionsChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsMemberSuggestionsChangePolicy">EventTypeArg.AsMemberSuggestionsChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsMicrosoftOfficeAddinChangePolicy">EventTypeArg.IsMicrosoftOfficeAddinChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsMicrosoftOfficeAddinChangePolicy">EventTypeArg.AsMicrosoftOfficeAddinChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsNetworkControlChangePolicy">EventTypeArg.IsNetworkControlChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsNetworkControlChangePolicy">EventTypeArg.AsNetworkControlChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperChangeDeploymentPolicy">EventTypeArg.IsPaperChangeDeploymentPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperChangeDeploymentPolicy">EventTypeArg.AsPaperChangeDeploymentPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperChangeMemberLinkPolicy">EventTypeArg.IsPaperChangeMemberLinkPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperChangeMemberLinkPolicy">EventTypeArg.AsPaperChangeMemberLinkPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperChangeMemberPolicy">EventTypeArg.IsPaperChangeMemberPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperChangeMemberPolicy">EventTypeArg.AsPaperChangeMemberPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperChangePolicy">EventTypeArg.IsPaperChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperChangePolicy">EventTypeArg.AsPaperChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperDefaultFolderPolicyChanged">EventTypeArg.IsPaperDefaultFolderPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperDefaultFolderPolicyChanged">EventTypeArg.AsPaperDefaultFolderPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperDesktopPolicyChanged">EventTypeArg.IsPaperDesktopPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperDesktopPolicyChanged">EventTypeArg.AsPaperDesktopPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperEnabledUsersGroupAddition">EventTypeArg.IsPaperEnabledUsersGroupAddition</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperEnabledUsersGroupAddition">EventTypeArg.AsPaperEnabledUsersGroupAddition</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPaperEnabledUsersGroupRemoval">EventTypeArg.IsPaperEnabledUsersGroupRemoval</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPaperEnabledUsersGroupRemoval">EventTypeArg.AsPaperEnabledUsersGroupRemoval</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPasswordStrengthRequirementsChangePolicy">EventTypeArg.IsPasswordStrengthRequirementsChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPasswordStrengthRequirementsChangePolicy">EventTypeArg.AsPasswordStrengthRequirementsChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsPermanentDeleteChangePolicy">EventTypeArg.IsPermanentDeleteChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsPermanentDeleteChangePolicy">EventTypeArg.AsPermanentDeleteChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsResellerSupportChangePolicy">EventTypeArg.IsResellerSupportChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsResellerSupportChangePolicy">EventTypeArg.AsResellerSupportChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsRewindPolicyChanged">EventTypeArg.IsRewindPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsRewindPolicyChanged">EventTypeArg.AsRewindPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSendForSignaturePolicyChanged">EventTypeArg.IsSendForSignaturePolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSendForSignaturePolicyChanged">EventTypeArg.AsSendForSignaturePolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharingChangeFolderJoinPolicy">EventTypeArg.IsSharingChangeFolderJoinPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharingChangeFolderJoinPolicy">EventTypeArg.AsSharingChangeFolderJoinPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharingChangeLinkAllowChangeExpirationPolicy">EventTypeArg.IsSharingChangeLinkAllowChangeExpirationPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharingChangeLinkAllowChangeExpirationPolicy">EventTypeArg.AsSharingChangeLinkAllowChangeExpirationPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharingChangeLinkDefaultExpirationPolicy">EventTypeArg.IsSharingChangeLinkDefaultExpirationPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharingChangeLinkDefaultExpirationPolicy">EventTypeArg.AsSharingChangeLinkDefaultExpirationPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharingChangeLinkEnforcePasswordPolicy">EventTypeArg.IsSharingChangeLinkEnforcePasswordPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharingChangeLinkEnforcePasswordPolicy">EventTypeArg.AsSharingChangeLinkEnforcePasswordPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharingChangeLinkPolicy">EventTypeArg.IsSharingChangeLinkPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharingChangeLinkPolicy">EventTypeArg.AsSharingChangeLinkPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSharingChangeMemberPolicy">EventTypeArg.IsSharingChangeMemberPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSharingChangeMemberPolicy">EventTypeArg.AsSharingChangeMemberPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsShowcaseChangeDownloadPolicy">EventTypeArg.IsShowcaseChangeDownloadPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsShowcaseChangeDownloadPolicy">EventTypeArg.AsShowcaseChangeDownloadPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsShowcaseChangeEnabledPolicy">EventTypeArg.IsShowcaseChangeEnabledPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsShowcaseChangeEnabledPolicy">EventTypeArg.AsShowcaseChangeEnabledPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsShowcaseChangeExternalSharingPolicy">EventTypeArg.IsShowcaseChangeExternalSharingPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsShowcaseChangeExternalSharingPolicy">EventTypeArg.AsShowcaseChangeExternalSharingPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSmarterSmartSyncPolicyChanged">EventTypeArg.IsSmarterSmartSyncPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSmarterSmartSyncPolicyChanged">EventTypeArg.AsSmarterSmartSyncPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSmartSyncChangePolicy">EventTypeArg.IsSmartSyncChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSmartSyncChangePolicy">EventTypeArg.AsSmartSyncChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSmartSyncNotOptOut">EventTypeArg.IsSmartSyncNotOptOut</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSmartSyncNotOptOut">EventTypeArg.AsSmartSyncNotOptOut</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSmartSyncOptOut">EventTypeArg.IsSmartSyncOptOut</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSmartSyncOptOut">EventTypeArg.AsSmartSyncOptOut</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsSsoChangePolicy">EventTypeArg.IsSsoChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsSsoChangePolicy">EventTypeArg.AsSsoChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamBrandingPolicyChanged">EventTypeArg.IsTeamBrandingPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamBrandingPolicyChanged">EventTypeArg.AsTeamBrandingPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamExtensionsPolicyChanged">EventTypeArg.IsTeamExtensionsPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamExtensionsPolicyChanged">EventTypeArg.AsTeamExtensionsPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamSelectiveSyncPolicyChanged">EventTypeArg.IsTeamSelectiveSyncPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamSelectiveSyncPolicyChanged">EventTypeArg.AsTeamSelectiveSyncPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamSharingWhitelistSubjectsChanged">EventTypeArg.IsTeamSharingWhitelistSubjectsChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamSharingWhitelistSubjectsChanged">EventTypeArg.AsTeamSharingWhitelistSubjectsChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTfaAddException">EventTypeArg.IsTfaAddException</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTfaAddException">EventTypeArg.AsTfaAddException</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTfaChangePolicy">EventTypeArg.IsTfaChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTfaChangePolicy">EventTypeArg.AsTfaChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTfaRemoveException">EventTypeArg.IsTfaRemoveException</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTfaRemoveException">EventTypeArg.AsTfaRemoveException</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTwoAccountChangePolicy">EventTypeArg.IsTwoAccountChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTwoAccountChangePolicy">EventTypeArg.AsTwoAccountChangePolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsViewerInfoPolicyChanged">EventTypeArg.IsViewerInfoPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsViewerInfoPolicyChanged">EventTypeArg.AsViewerInfoPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsWatermarkingPolicyChanged">EventTypeArg.IsWatermarkingPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsWatermarkingPolicyChanged">EventTypeArg.AsWatermarkingPolicyChanged</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsWebSessionsChangeActiveSessionLimit">EventTypeArg.IsWebSessionsChangeActiveSessionLimit</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsWebSessionsChangeActiveSessionLimit">EventTypeArg.AsWebSessionsChangeActiveSessionLimit</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsWebSessionsChangeFixedLengthPolicy">EventTypeArg.IsWebSessionsChangeFixedLengthPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsWebSessionsChangeFixedLengthPolicy">EventTypeArg.AsWebSessionsChangeFixedLengthPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsWebSessionsChangeIdleLengthPolicy">EventTypeArg.IsWebSessionsChangeIdleLengthPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsWebSessionsChangeIdleLengthPolicy">EventTypeArg.AsWebSessionsChangeIdleLengthPolicy</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDataResidencyMigrationRequestSuccessful">EventTypeArg.IsDataResidencyMigrationRequestSuccessful</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDataResidencyMigrationRequestSuccessful">EventTypeArg.AsDataResidencyMigrationRequestSuccessful</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsDataResidencyMigrationRequestUnsuccessful">EventTypeArg.IsDataResidencyMigrationRequestUnsuccessful</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsDataResidencyMigrationRequestUnsuccessful">EventTypeArg.AsDataResidencyMigrationRequestUnsuccessful</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamMergeFrom">EventTypeArg.IsTeamMergeFrom</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamMergeFrom">EventTypeArg.AsTeamMergeFrom</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamMergeTo">EventTypeArg.IsTeamMergeTo</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamMergeTo">EventTypeArg.AsTeamMergeTo</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamProfileAddBackground">EventTypeArg.IsTeamProfileAddBackground</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamProfileAddBackground">EventTypeArg.AsTeamProfileAddBackground</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamProfileAddLogo">EventTypeArg.IsTeamProfileAddLogo</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamProfileAddLogo">EventTypeArg.AsTeamProfileAddLogo</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamProfileChangeBackground">EventTypeArg.IsTeamProfileChangeBackground</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamProfileChangeBackground">EventTypeArg.AsTeamProfileChangeBackground</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamProfileChangeDefaultLanguage">EventTypeArg.IsTeamProfileChangeDefaultLanguage</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamProfileChangeDefaultLanguage">EventTypeArg.AsTeamProfileChangeDefaultLanguage</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamProfileChangeLogo">EventTypeArg.IsTeamProfileChangeLogo</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamProfileChangeLogo">EventTypeArg.AsTeamProfileChangeLogo</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamProfileChangeName">EventTypeArg.IsTeamProfileChangeName</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamProfileChangeName">EventTypeArg.AsTeamProfileChangeName</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamProfileRemoveBackground">EventTypeArg.IsTeamProfileRemoveBackground</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamProfileRemoveBackground">EventTypeArg.AsTeamProfileRemoveBackground</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamProfileRemoveLogo">EventTypeArg.IsTeamProfileRemoveLogo</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamProfileRemoveLogo">EventTypeArg.AsTeamProfileRemoveLogo</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTfaAddBackupPhone">EventTypeArg.IsTfaAddBackupPhone</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTfaAddBackupPhone">EventTypeArg.AsTfaAddBackupPhone</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTfaAddSecurityKey">EventTypeArg.IsTfaAddSecurityKey</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTfaAddSecurityKey">EventTypeArg.AsTfaAddSecurityKey</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTfaChangeBackupPhone">EventTypeArg.IsTfaChangeBackupPhone</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTfaChangeBackupPhone">EventTypeArg.AsTfaChangeBackupPhone</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTfaChangeStatus">EventTypeArg.IsTfaChangeStatus</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTfaChangeStatus">EventTypeArg.AsTfaChangeStatus</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTfaRemoveBackupPhone">EventTypeArg.IsTfaRemoveBackupPhone</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTfaRemoveBackupPhone">EventTypeArg.AsTfaRemoveBackupPhone</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTfaRemoveSecurityKey">EventTypeArg.IsTfaRemoveSecurityKey</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTfaRemoveSecurityKey">EventTypeArg.AsTfaRemoveSecurityKey</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTfaReset">EventTypeArg.IsTfaReset</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTfaReset">EventTypeArg.AsTfaReset</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsChangedEnterpriseAdminRole">EventTypeArg.IsChangedEnterpriseAdminRole</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsChangedEnterpriseAdminRole">EventTypeArg.AsChangedEnterpriseAdminRole</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsChangedEnterpriseConnectedTeamStatus">EventTypeArg.IsChangedEnterpriseConnectedTeamStatus</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsChangedEnterpriseConnectedTeamStatus">EventTypeArg.AsChangedEnterpriseConnectedTeamStatus</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsEndedEnterpriseAdminSession">EventTypeArg.IsEndedEnterpriseAdminSession</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsEndedEnterpriseAdminSession">EventTypeArg.AsEndedEnterpriseAdminSession</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsEndedEnterpriseAdminSessionDeprecated">EventTypeArg.IsEndedEnterpriseAdminSessionDeprecated</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsEndedEnterpriseAdminSessionDeprecated">EventTypeArg.AsEndedEnterpriseAdminSessionDeprecated</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsEnterpriseSettingsLocking">EventTypeArg.IsEnterpriseSettingsLocking</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsEnterpriseSettingsLocking">EventTypeArg.AsEnterpriseSettingsLocking</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsGuestAdminChangeStatus">EventTypeArg.IsGuestAdminChangeStatus</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsGuestAdminChangeStatus">EventTypeArg.AsGuestAdminChangeStatus</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsStartedEnterpriseAdminSession">EventTypeArg.IsStartedEnterpriseAdminSession</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsStartedEnterpriseAdminSession">EventTypeArg.AsStartedEnterpriseAdminSession</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamMergeRequestAccepted">EventTypeArg.IsTeamMergeRequestAccepted</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamMergeRequestAccepted">EventTypeArg.AsTeamMergeRequestAccepted</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamMergeRequestAcceptedShownToPrimaryTeam">EventTypeArg.IsTeamMergeRequestAcceptedShownToPrimaryTeam</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamMergeRequestAcceptedShownToPrimaryTeam">EventTypeArg.AsTeamMergeRequestAcceptedShownToPrimaryTeam</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamMergeRequestAcceptedShownToSecondaryTeam">EventTypeArg.IsTeamMergeRequestAcceptedShownToSecondaryTeam</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamMergeRequestAcceptedShownToSecondaryTeam">EventTypeArg.AsTeamMergeRequestAcceptedShownToSecondaryTeam</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamMergeRequestAutoCanceled">EventTypeArg.IsTeamMergeRequestAutoCanceled</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamMergeRequestAutoCanceled">EventTypeArg.AsTeamMergeRequestAutoCanceled</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamMergeRequestCanceled">EventTypeArg.IsTeamMergeRequestCanceled</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamMergeRequestCanceled">EventTypeArg.AsTeamMergeRequestCanceled</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamMergeRequestCanceledShownToPrimaryTeam">EventTypeArg.IsTeamMergeRequestCanceledShownToPrimaryTeam</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamMergeRequestCanceledShownToPrimaryTeam">EventTypeArg.AsTeamMergeRequestCanceledShownToPrimaryTeam</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamMergeRequestCanceledShownToSecondaryTeam">EventTypeArg.IsTeamMergeRequestCanceledShownToSecondaryTeam</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamMergeRequestCanceledShownToSecondaryTeam">EventTypeArg.AsTeamMergeRequestCanceledShownToSecondaryTeam</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamMergeRequestExpired">EventTypeArg.IsTeamMergeRequestExpired</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamMergeRequestExpired">EventTypeArg.AsTeamMergeRequestExpired</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamMergeRequestExpiredShownToPrimaryTeam">EventTypeArg.IsTeamMergeRequestExpiredShownToPrimaryTeam</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamMergeRequestExpiredShownToPrimaryTeam">EventTypeArg.AsTeamMergeRequestExpiredShownToPrimaryTeam</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamMergeRequestExpiredShownToSecondaryTeam">EventTypeArg.IsTeamMergeRequestExpiredShownToSecondaryTeam</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamMergeRequestExpiredShownToSecondaryTeam">EventTypeArg.AsTeamMergeRequestExpiredShownToSecondaryTeam</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamMergeRequestRejectedShownToPrimaryTeam">EventTypeArg.IsTeamMergeRequestRejectedShownToPrimaryTeam</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamMergeRequestRejectedShownToPrimaryTeam">EventTypeArg.AsTeamMergeRequestRejectedShownToPrimaryTeam</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamMergeRequestRejectedShownToSecondaryTeam">EventTypeArg.IsTeamMergeRequestRejectedShownToSecondaryTeam</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamMergeRequestRejectedShownToSecondaryTeam">EventTypeArg.AsTeamMergeRequestRejectedShownToSecondaryTeam</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamMergeRequestReminder">EventTypeArg.IsTeamMergeRequestReminder</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamMergeRequestReminder">EventTypeArg.AsTeamMergeRequestReminder</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamMergeRequestReminderShownToPrimaryTeam">EventTypeArg.IsTeamMergeRequestReminderShownToPrimaryTeam</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamMergeRequestReminderShownToPrimaryTeam">EventTypeArg.AsTeamMergeRequestReminderShownToPrimaryTeam</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamMergeRequestReminderShownToSecondaryTeam">EventTypeArg.IsTeamMergeRequestReminderShownToSecondaryTeam</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamMergeRequestReminderShownToSecondaryTeam">EventTypeArg.AsTeamMergeRequestReminderShownToSecondaryTeam</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamMergeRequestRevoked">EventTypeArg.IsTeamMergeRequestRevoked</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamMergeRequestRevoked">EventTypeArg.AsTeamMergeRequestRevoked</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamMergeRequestSentShownToPrimaryTeam">EventTypeArg.IsTeamMergeRequestSentShownToPrimaryTeam</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamMergeRequestSentShownToPrimaryTeam">EventTypeArg.AsTeamMergeRequestSentShownToPrimaryTeam</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsTeamMergeRequestSentShownToSecondaryTeam">EventTypeArg.IsTeamMergeRequestSentShownToSecondaryTeam</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsTeamMergeRequestSentShownToSecondaryTeam">EventTypeArg.AsTeamMergeRequestSentShownToSecondaryTeam</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_IsOther">EventTypeArg.IsOther</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.html#Dropbox_Api_TeamLog_EventTypeArg_AsOther">EventTypeArg.AsOther</a>
    </div>
    <div>
      <span class="xref">System.Object.Equals(System.Object)</span>
    </div>
    <div>
      <span class="xref">System.Object.Equals(System.Object, System.Object)</span>
    </div>
    <div>
      <span class="xref">System.Object.GetHashCode()</span>
    </div>
    <div>
      <span class="xref">System.Object.GetType()</span>
    </div>
    <div>
      <span class="xref">System.Object.MemberwiseClone()</span>
    </div>
    <div>
      <span class="xref">System.Object.ReferenceEquals(System.Object, System.Object)</span>
    </div>
    <div>
      <span class="xref">System.Object.ToString()</span>
    </div>
  </div>
  <h6><strong>Namespace</strong>: <a class="xref" href="Dropbox.Api.TeamLog.html">Dropbox.Api.TeamLog</a></h6>
  <h6><strong>Assembly</strong>: Dropbox.Api.dll</h6>
  <h5 id="Dropbox_Api_TeamLog_EventTypeArg_SharedLinkRemoveExpiry_syntax">Syntax</h5>
  <div class="codewrapper">
    <pre><code class="lang-csharp hljs">public sealed class SharedLinkRemoveExpiry : EventTypeArg</code></pre>
  </div>
  <h3 id="fields">Fields
  </h3>
  <span class="small pull-right mobile-hide">
    <span class="divider">|</span>
    <a href="https://github.com/dropbox/dropbox-sdk-dotnet/new/doc_fx_integration/apiSpec/new?filename=Dropbox_Api_TeamLog_EventTypeArg_SharedLinkRemoveExpiry_Instance.md&amp;value=---%0Auid%3A%20Dropbox.Api.TeamLog.EventTypeArg.SharedLinkRemoveExpiry.Instance%0Asummary%3A%20'*You%20can%20override%20summary%20for%20the%20API%20here%20using%20*MARKDOWN*%20syntax'%0A---%0A%0A*Please%20type%20below%20more%20information%20about%20this%20API%3A*%0A%0A">Improve this Doc</a>
  </span>
  <span class="small pull-right mobile-hide">
    <a href="https://github.com/dropbox/dropbox-sdk-dotnet/blob/doc_fx_integration/dropbox-sdk-dotnet/Dropbox.Api/Generated/TeamLog/EventTypeArg.cs/#L35939">View Source</a>
  </span>
  <h4 id="Dropbox_Api_TeamLog_EventTypeArg_SharedLinkRemoveExpiry_Instance" data-uid="Dropbox.Api.TeamLog.EventTypeArg.SharedLinkRemoveExpiry.Instance">Instance</h4>
  <div class="markdown level1 summary"><p>A singleton instance of SharedLinkRemoveExpiry</p>
</div>
  <div class="markdown level1 conceptual"></div>
  <h5 class="decalaration">Declaration</h5>
  <div class="codewrapper">
    <pre><code class="lang-csharp hljs">public static readonly EventTypeArg.SharedLinkRemoveExpiry Instance</code></pre>
  </div>
  <h5 class="fieldValue">Field Value</h5>
  <table class="table table-bordered table-striped table-condensed">
    <thead>
      <tr>
        <th>Type</th>
        <th>Description</th>
      </tr>
    </thead>
    <tbody>
      <tr>
        <td><a class="xref" href="Dropbox.Api.TeamLog.EventTypeArg.SharedLinkRemoveExpiry.html">EventTypeArg.SharedLinkRemoveExpiry</a></td>
        <td></td>
      </tr>
    </tbody>
  </table>
</article>
          </div>
          
          <div class="hidden-sm col-md-2" role="complementary">
            <div class="sideaffix">
              <div class="contribution">
                <ul class="nav">
                  <li>
                    <a href="https://github.com/dropbox/dropbox-sdk-dotnet/new/doc_fx_integration/apiSpec/new?filename=Dropbox_Api_TeamLog_EventTypeArg_SharedLinkRemoveExpiry.md&amp;value=---%0Auid%3A%20Dropbox.Api.TeamLog.EventTypeArg.SharedLinkRemoveExpiry%0Asummary%3A%20'*You%20can%20override%20summary%20for%20the%20API%20here%20using%20*MARKDOWN*%20syntax'%0A---%0A%0A*Please%20type%20below%20more%20information%20about%20this%20API%3A*%0A%0A" class="contribution-link">Improve this Doc</a>
                  </li>
                  <li>
                    <a href="https://github.com/dropbox/dropbox-sdk-dotnet/blob/doc_fx_integration/dropbox-sdk-dotnet/Dropbox.Api/Generated/TeamLog/EventTypeArg.cs/#L35914" class="contribution-link">View Source</a>
                  </li>
                </ul>
              </div>
              <nav class="bs-docs-sidebar hidden-print hidden-xs hidden-sm affix" id="affix">
                <h5>In This Article</h5>
                <div></div>
              </nav>
            </div>
          </div>
        </div>
      </div>
      
      <footer>
        <div class="grad-bottom"></div>
        <div class="footer">
          <div class="container">
            <span class="pull-right">
              <a href="#top">Back to top</a>
            </span>
            
            <span>Generated by <strong>DocFX</strong></span>
          </div>
        </div>
      </footer>
    </div>
    
    <script type="text/javascript" src="../../../styles/docfx.vendor.js"></script>
    <script type="text/javascript" src="../../../styles/docfx.js"></script>
    <script type="text/javascript" src="../../../styles/main.js"></script>
  </body>
</html>
