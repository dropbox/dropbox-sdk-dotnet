<!DOCTYPE html>
<!--[if IE]><![endif]-->
<html>
  
  <head>
    <meta charset="utf-8">
    <meta http-equiv="X-UA-Compatible" content="IE=edge,chrome=1">
    <title>Class FileLockingPolicyState.Enabled
   </title>
    <meta name="viewport" content="width=device-width">
    <meta name="title" content="Class FileLockingPolicyState.Enabled
   ">
    <meta name="generator" content="docfx 2.58.4.0">
    
    <link rel="shortcut icon" href="../../../favicon.ico">
    <link rel="stylesheet" href="../../../styles/docfx.vendor.css">
    <link rel="stylesheet" href="../../../styles/docfx.css">
    <link rel="stylesheet" href="../../../styles/main.css">
    <meta property="docfx:navrel" content="../../../toc.html">
    <meta property="docfx:tocrel" content="toc.html">
    
    
    
  </head>
  <body data-spy="scroll" data-target="#affix" data-offset="120">
    <div id="wrapper">
      <header>
        
        <nav id="autocollapse" class="navbar navbar-inverse ng-scope" role="navigation">
          <div class="container">
            <div class="navbar-header">
              <button type="button" class="navbar-toggle" data-toggle="collapse" data-target="#navbar">
                <span class="sr-only">Toggle navigation</span>
                <span class="icon-bar"></span>
                <span class="icon-bar"></span>
                <span class="icon-bar"></span>
              </button>
              
              <a class="navbar-brand" href="../../../index.html">
                <img id="logo" class="svg" src="../../../logo.svg" alt="">
              </a>
            </div>
            <div class="collapse navbar-collapse" id="navbar">
              <form class="navbar-form navbar-right" role="search" id="search">
                <div class="form-group">
                  <input type="text" class="form-control" id="search-query" placeholder="Search" autocomplete="off">
                </div>
              </form>
            </div>
          </div>
        </nav>
        
        <div class="subnav navbar navbar-default">
          <div class="container hide-when-search" id="breadcrumb">
            <ul class="breadcrumb">
              <li></li>
            </ul>
          </div>
        </div>
      </header>
      <div role="main" class="container body-content hide-when-search">
        
        <div class="sidenav hide-when-search">
          <a class="btn toc-toggle collapse" data-toggle="collapse" href="#sidetoggle" aria-expanded="false" aria-controls="sidetoggle">Show / Hide Table of Contents</a>
          <div class="sidetoggle collapse" id="sidetoggle">
            <div id="sidetoc"></div>
          </div>
        </div>
        <div class="article row grid-right">
          <div class="col-md-10">
            <article class="content wrap" id="_content" data-uid="Dropbox.Api.TeamPolicies.FileLockingPolicyState.Enabled">
  
  
  <h1 id="Dropbox_Api_TeamPolicies_FileLockingPolicyState_Enabled" data-uid="Dropbox.Api.TeamPolicies.FileLockingPolicyState.Enabled" class="text-break">Class FileLockingPolicyState.Enabled
  </h1>
  <div class="markdown level0 summary"><p>File locking feature is allowed.</p>
</div>
  <div class="markdown level0 conceptual"></div>
  <div class="inheritance">
    <h5>Inheritance</h5>
    <div class="level0"><span class="xref">System.Object</span></div>
    <div class="level1"><a class="xref" href="Dropbox.Api.TeamPolicies.FileLockingPolicyState.html">FileLockingPolicyState</a></div>
    <div class="level2"><span class="xref">FileLockingPolicyState.Enabled</span></div>
  </div>
  <div class="inheritedMembers">
    <h5>Inherited Members</h5>
    <div>
      <a class="xref" href="Dropbox.Api.TeamPolicies.FileLockingPolicyState.html#Dropbox_Api_TeamPolicies_FileLockingPolicyState_IsDisabled">FileLockingPolicyState.IsDisabled</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamPolicies.FileLockingPolicyState.html#Dropbox_Api_TeamPolicies_FileLockingPolicyState_AsDisabled">FileLockingPolicyState.AsDisabled</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamPolicies.FileLockingPolicyState.html#Dropbox_Api_TeamPolicies_FileLockingPolicyState_IsEnabled">FileLockingPolicyState.IsEnabled</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamPolicies.FileLockingPolicyState.html#Dropbox_Api_TeamPolicies_FileLockingPolicyState_AsEnabled">FileLockingPolicyState.AsEnabled</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamPolicies.FileLockingPolicyState.html#Dropbox_Api_TeamPolicies_FileLockingPolicyState_IsOther">FileLockingPolicyState.IsOther</a>
    </div>
    <div>
      <a class="xref" href="Dropbox.Api.TeamPolicies.FileLockingPolicyState.html#Dropbox_Api_TeamPolicies_FileLockingPolicyState_AsOther">FileLockingPolicyState.AsOther</a>
    </div>
    <div>
      <span class="xref">System.Object.Equals(System.Object)</span>
    </div>
    <div>
      <span class="xref">System.Object.Equals(System.Object, System.Object)</span>
    </div>
    <div>
      <span class="xref">System.Object.GetHashCode()</span>
    </div>
    <div>
      <span class="xref">System.Object.GetType()</span>
    </div>
    <div>
      <span class="xref">System.Object.MemberwiseClone()</span>
    </div>
    <div>
      <span class="xref">System.Object.ReferenceEquals(System.Object, System.Object)</span>
    </div>
    <div>
      <span class="xref">System.Object.ToString()</span>
    </div>
  </div>
  <h6><strong>Namespace</strong>: <a class="xref" href="Dropbox.Api.TeamPolicies.html">Dropbox.Api.TeamPolicies</a></h6>
  <h6><strong>Assembly</strong>: Dropbox.Api.dll</h6>
  <h5 id="Dropbox_Api_TeamPolicies_FileLockingPolicyState_Enabled_syntax">Syntax</h5>
  <div class="codewrapper">
    <pre><code class="lang-csharp hljs">public sealed class Enabled : FileLockingPolicyState</code></pre>
  </div>
  <h3 id="fields">Fields
  </h3>
  <span class="small pull-right mobile-hide">
    <span class="divider">|</span>
    <a href="https://github.com/dropbox/dropbox-sdk-dotnet/new/doc_fx_integration/apiSpec/new?filename=Dropbox_Api_TeamPolicies_FileLockingPolicyState_Enabled_Instance.md&amp;value=---%0Auid%3A%20Dropbox.Api.TeamPolicies.FileLockingPolicyState.Enabled.Instance%0Asummary%3A%20'*You%20can%20override%20summary%20for%20the%20API%20here%20using%20*MARKDOWN*%20syntax'%0A---%0A%0A*Please%20type%20below%20more%20information%20about%20this%20API%3A*%0A%0A">Improve this Doc</a>
  </span>
  <span class="small pull-right mobile-hide">
    <a href="https://github.com/dropbox/dropbox-sdk-dotnet/blob/doc_fx_integration/dropbox-sdk-dotnet/Dropbox.Api/Generated/TeamPolicies/FileLockingPolicyState.cs/#L277">View Source</a>
  </span>
  <h4 id="Dropbox_Api_TeamPolicies_FileLockingPolicyState_Enabled_Instance" data-uid="Dropbox.Api.TeamPolicies.FileLockingPolicyState.Enabled.Instance">Instance</h4>
  <div class="markdown level1 summary"><p>A singleton instance of Enabled</p>
</div>
  <div class="markdown level1 conceptual"></div>
  <h5 class="decalaration">Declaration</h5>
  <div class="codewrapper">
    <pre><code class="lang-csharp hljs">public static readonly FileLockingPolicyState.Enabled Instance</code></pre>
  </div>
  <h5 class="fieldValue">Field Value</h5>
  <table class="table table-bordered table-striped table-condensed">
    <thead>
      <tr>
        <th>Type</th>
        <th>Description</th>
      </tr>
    </thead>
    <tbody>
      <tr>
        <td><a class="xref" href="Dropbox.Api.TeamPolicies.FileLockingPolicyState.Enabled.html">FileLockingPolicyState.Enabled</a></td>
        <td></td>
      </tr>
    </tbody>
  </table>
</article>
          </div>
          
          <div class="hidden-sm col-md-2" role="complementary">
            <div class="sideaffix">
              <div class="contribution">
                <ul class="nav">
                  <li>
                    <a href="https://github.com/dropbox/dropbox-sdk-dotnet/new/doc_fx_integration/apiSpec/new?filename=Dropbox_Api_TeamPolicies_FileLockingPolicyState_Enabled.md&amp;value=---%0Auid%3A%20Dropbox.Api.TeamPolicies.FileLockingPolicyState.Enabled%0Asummary%3A%20'*You%20can%20override%20summary%20for%20the%20API%20here%20using%20*MARKDOWN*%20syntax'%0A---%0A%0A*Please%20type%20below%20more%20information%20about%20this%20API%3A*%0A%0A" class="contribution-link">Improve this Doc</a>
                  </li>
                  <li>
                    <a href="https://github.com/dropbox/dropbox-sdk-dotnet/blob/doc_fx_integration/dropbox-sdk-dotnet/Dropbox.Api/Generated/TeamPolicies/FileLockingPolicyState.cs/#L253" class="contribution-link">View Source</a>
                  </li>
                </ul>
              </div>
              <nav class="bs-docs-sidebar hidden-print hidden-xs hidden-sm affix" id="affix">
                <h5>In This Article</h5>
                <div></div>
              </nav>
            </div>
          </div>
        </div>
      </div>
      
      <footer>
        <div class="grad-bottom"></div>
        <div class="footer">
          <div class="container">
            <span class="pull-right">
              <a href="#top">Back to top</a>
            </span>
            
            <span>Generated by <strong>DocFX</strong></span>
          </div>
        </div>
      </footer>
    </div>
    
    <script type="text/javascript" src="../../../styles/docfx.vendor.js"></script>
    <script type="text/javascript" src="../../../styles/docfx.js"></script>
    <script type="text/javascript" src="../../../styles/main.js"></script>
  </body>
</html>
